library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_char_l is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(11 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_char_l is
	type rom is array(0 to  4095) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",X"00",X"18",X"1C",X"18",X"18",X"18",X"18",X"3C",
		X"00",X"7C",X"E6",X"C6",X"30",X"0C",X"C6",X"7E",X"00",X"7C",X"C6",X"C0",X"70",X"C6",X"C6",X"7C",
		X"00",X"68",X"68",X"6C",X"64",X"FE",X"60",X"F0",X"00",X"7E",X"02",X"7E",X"C2",X"C0",X"C6",X"7C",
		X"00",X"7C",X"C6",X"06",X"7E",X"C6",X"C6",X"7C",X"00",X"FE",X"C2",X"C2",X"60",X"30",X"18",X"18",
		X"00",X"7C",X"C6",X"C6",X"7C",X"C6",X"C6",X"7C",X"00",X"7C",X"C6",X"C6",X"FC",X"C0",X"C6",X"7C",
		X"00",X"70",X"58",X"C8",X"CC",X"FC",X"C6",X"C6",X"00",X"7E",X"CC",X"CC",X"7C",X"CC",X"CC",X"7E",
		X"00",X"78",X"CC",X"06",X"06",X"86",X"CC",X"78",X"00",X"3E",X"6C",X"CC",X"CC",X"CC",X"6C",X"3E",
		X"00",X"FE",X"CC",X"0C",X"3C",X"0C",X"CC",X"FE",X"00",X"FE",X"CC",X"0C",X"3C",X"0C",X"0C",X"1E",
		X"00",X"78",X"CC",X"06",X"06",X"E6",X"CC",X"78",X"00",X"EE",X"6C",X"6C",X"7C",X"6C",X"6C",X"EE",
		X"00",X"3C",X"18",X"18",X"18",X"18",X"18",X"3C",X"00",X"F0",X"60",X"60",X"60",X"60",X"6C",X"38",
		X"00",X"9E",X"CC",X"6C",X"3C",X"6C",X"CC",X"DE",X"00",X"1E",X"0C",X"0C",X"0C",X"0C",X"CC",X"FE",
		X"00",X"C6",X"EE",X"FE",X"D6",X"D6",X"C6",X"C6",X"00",X"C6",X"CE",X"DE",X"F6",X"E6",X"C6",X"C6",
		X"00",X"7C",X"C6",X"C6",X"C6",X"C6",X"C6",X"7C",X"00",X"7E",X"CC",X"CC",X"7C",X"0C",X"0C",X"1E",
		X"00",X"38",X"6C",X"C6",X"C6",X"D6",X"6C",X"D8",X"00",X"7E",X"CC",X"CC",X"7C",X"6C",X"CC",X"DE",
		X"00",X"7C",X"8E",X"1C",X"78",X"F0",X"E2",X"7C",X"00",X"7E",X"5A",X"18",X"18",X"18",X"18",X"3C",
		X"00",X"DE",X"8C",X"8C",X"8C",X"8C",X"8C",X"78",X"00",X"DE",X"8C",X"8C",X"8C",X"58",X"58",X"30",
		X"00",X"B6",X"B6",X"B6",X"B6",X"FE",X"6C",X"28",X"00",X"C6",X"6E",X"3C",X"38",X"78",X"EC",X"C6",
		X"00",X"E6",X"6C",X"78",X"30",X"30",X"18",X"1C",X"00",X"FE",X"E6",X"70",X"38",X"1C",X"CE",X"FE",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"10",X"00",X"00",X"00",
		X"00",X"00",X"10",X"00",X"00",X"10",X"00",X"00",X"00",X"0C",X"12",X"14",X"08",X"14",X"22",X"7C",
		X"30",X"30",X"38",X"38",X"18",X"08",X"00",X"04",X"38",X"44",X"44",X"20",X"10",X"10",X"00",X"10",
		X"00",X"20",X"10",X"08",X"08",X"08",X"10",X"20",X"00",X"08",X"10",X"20",X"20",X"20",X"10",X"08",
		X"00",X"10",X"10",X"10",X"FE",X"10",X"10",X"10",X"00",X"00",X"00",X"00",X"7E",X"00",X"00",X"00",
		X"00",X"00",X"7E",X"00",X"00",X"7E",X"00",X"00",X"00",X"44",X"EE",X"EE",X"FE",X"7C",X"38",X"10",
		X"38",X"44",X"44",X"38",X"10",X"7C",X"10",X"10",X"10",X"38",X"54",X"10",X"38",X"44",X"44",X"38",
		X"18",X"38",X"28",X"48",X"28",X"0C",X"0E",X"06",X"10",X"38",X"7C",X"54",X"FE",X"28",X"44",X"28",
		X"00",X"00",X"A7",X"A9",X"A7",X"A5",X"49",X"00",X"00",X"00",X"02",X"06",X"0A",X"0A",X"06",X"00",
		X"00",X"00",X"07",X"31",X"53",X"51",X"57",X"00",X"00",X"04",X"04",X"06",X"05",X"05",X"06",X"00",
		X"00",X"00",X"00",X"FF",X"FF",X"00",X"00",X"00",X"10",X"38",X"7C",X"FE",X"38",X"38",X"38",X"38",
		X"3C",X"42",X"99",X"85",X"85",X"99",X"42",X"3C",X"00",X"7C",X"18",X"F0",X"FC",X"00",X"00",X"00",
		X"00",X"00",X"00",X"01",X"0F",X"7F",X"00",X"00",X"00",X"3E",X"0C",X"F8",X"FE",X"80",X"00",X"00",
		X"00",X"00",X"00",X"00",X"07",X"3F",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"03",X"02",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"02",
		X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"02",X"02",X"02",X"02",X"02",X"02",X"02",X"03",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"40",X"00",X"20",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"10",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"08",
		X"00",X"00",X"00",X"00",X"00",X"04",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",
		X"00",X"00",X"00",X"08",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"80",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"80",X"80",X"80",X"80",X"80",X"80",X"80",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"00",X"00",X"C8",X"C8",X"C8",X"C8",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"20",X"20",X"30",X"31",X"FD",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"79",X"79",X"79",X"79",X"00",X"00",X"3E",X"7C",X"78",X"F8",X"F0",X"F0",X"F0",X"F0",
		X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"E0",X"00",X"00",X"18",X"18",X"18",X"18",X"3C",X"3C",
		X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"FF",X"FF",X"00",X"00",X"7E",X"7E",X"7E",X"7E",X"00",X"00",
		X"00",X"00",X"3C",X"00",X"3C",X"3C",X"00",X"00",X"3C",X"00",X"00",X"3C",X"3C",X"00",X"00",X"3C",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"04",X"04",X"0C",X"8C",X"BE",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"9E",X"9E",X"9E",X"9E",X"00",X"00",X"7C",X"3E",X"1E",X"1F",X"0F",X"0F",X"0F",X"0F",
		X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"07",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"00",X"00",X"13",X"13",X"13",X"13",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"7E",X"7E",X"FF",X"7E",X"7E",X"FF",X"7E",X"7E",
		X"C0",X"60",X"F0",X"78",X"7C",X"FE",X"7F",X"7E",X"03",X"06",X"0F",X"1E",X"3E",X"7F",X"FE",X"7E",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"C0",X"70",X"FC",X"7F",X"7F",X"FF",X"7F",X"7F",
		X"03",X"0E",X"3F",X"FE",X"FE",X"FF",X"FE",X"FE",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",
		X"FF",X"FF",X"CC",X"CC",X"CC",X"CC",X"FF",X"FF",X"00",X"80",X"40",X"20",X"10",X"88",X"C4",X"F2",
		X"F1",X"E8",X"E8",X"D0",X"A3",X"47",X"8F",X"1F",X"FF",X"00",X"00",X"F0",X"E3",X"C7",X"8F",X"1F",
		X"2F",X"2F",X"17",X"8B",X"C5",X"E2",X"F1",X"F8",X"FF",X"00",X"00",X"0F",X"C7",X"E3",X"F1",X"F8",
		X"74",X"74",X"F8",X"D0",X"A3",X"47",X"8F",X"1F",X"00",X"01",X"02",X"04",X"08",X"11",X"23",X"47",
		X"8F",X"17",X"17",X"0B",X"C5",X"E2",X"F1",X"F8",X"00",X"00",X"80",X"C0",X"E0",X"70",X"38",X"1C",
		X"1C",X"8E",X"AE",X"FE",X"DE",X"DF",X"FF",X"FF",X"07",X"07",X"07",X"06",X"0E",X"0E",X"0E",X"1C",
		X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"E0",X"F8",X"3C",X"1C",X"0C",X"0C",X"0C",
		X"E0",X"FE",X"FF",X"07",X"41",X"E0",X"A8",X"BC",X"F5",X"F7",X"BE",X"BE",X"F7",X"F7",X"BE",X"BE",
		X"00",X"00",X"CE",X"CE",X"CE",X"C0",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"3E",X"1C",X"1C",X"1C",X"07",X"7F",X"FF",X"E0",X"82",X"07",X"15",X"3D",
		X"AF",X"EF",X"7D",X"7D",X"EF",X"EF",X"7D",X"7D",X"00",X"00",X"73",X"73",X"73",X"03",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"7C",X"38",X"38",X"38",
		X"00",X"00",X"01",X"03",X"07",X"0E",X"1C",X"38",X"38",X"71",X"75",X"7F",X"7B",X"FB",X"FF",X"FF",
		X"E0",X"E0",X"E0",X"60",X"70",X"70",X"70",X"38",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",
		X"03",X"07",X"1F",X"3C",X"38",X"30",X"30",X"30",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"80",X"80",X"80",
		X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"F0",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"01",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",X"0F",
		X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"3E",X"1C",X"7E",X"7E",X"FF",X"7E",X"7E",X"FF",X"7E",X"7E",
		X"C0",X"60",X"F0",X"78",X"7C",X"FE",X"7F",X"7E",X"03",X"09",X"0F",X"1E",X"3E",X"7F",X"FE",X"7E",
		X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"C0",X"70",X"FC",X"7F",X"7F",X"FF",X"7F",X"7F",
		X"03",X"0E",X"3F",X"FE",X"FE",X"FF",X"FE",X"FE",X"00",X"00",X"00",X"00",X"03",X"0F",X"3F",X"FF",
		X"00",X"00",X"80",X"C5",X"C7",X"05",X"10",X"71",X"00",X"00",X"00",X"80",X"C0",X"C0",X"10",X"10",
		X"00",X"00",X"00",X"01",X"03",X"03",X"02",X"18",X"00",X"00",X"00",X"00",X"00",X"00",X"C0",X"10",
		X"00",X"00",X"00",X"00",X"60",X"70",X"01",X"70",X"00",X"00",X"01",X"03",X"07",X"00",X"80",X"38",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"00",X"C0",X"F0",X"F8",X"FC",X"FE",X"FE",X"FF",
		X"C0",X"E9",X"E5",X"F4",X"72",X"79",X"38",X"3C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"F8",X"FC",X"FE",X"7F",X"7C",X"F8",X"E0",X"E0",
		X"7E",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"81",X"81",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"81",X"00",X"00",X"00",X"00",X"C3",X"FF",X"00",X"03",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",
		X"01",X"53",X"13",X"27",X"26",X"4E",X"0C",X"1C",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"1F",X"3F",X"7F",X"FF",X"3F",X"1F",X"07",X"07",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",
		X"81",X"DB",X"7E",X"24",X"24",X"7E",X"E7",X"C3",X"80",X"D8",X"70",X"32",X"3E",X"7C",X"E6",X"C3",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"4E",X"FF",X"00",X"00",X"00",X"80",X"80",X"C0",X"E0",X"F0",
		X"FF",X"FF",X"0F",X"EE",X"EE",X"DE",X"DC",X"BC",X"B8",X"78",X"70",X"F0",X"E0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"F0",X"90",X"98",X"88",X"CC",X"44",X"46",X"63",X"21",X"30",X"18",X"0C",X"FF",
		X"FF",X"FF",X"F8",X"FB",X"FB",X"F7",X"F7",X"F7",X"EF",X"EF",X"E0",X"FF",X"FF",X"F7",X"F7",X"F7",
		X"11",X"11",X"11",X"22",X"22",X"24",X"24",X"24",X"24",X"24",X"FF",X"FF",X"FF",X"FF",X"24",X"24",
		X"00",X"00",X"00",X"FF",X"99",X"99",X"18",X"18",X"18",X"3C",X"3C",X"3C",X"3C",X"7E",X"7E",X"FF",
		X"FF",X"FF",X"00",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"7E",X"00",X"FF",X"FF",X"7E",X"7E",X"7E",
		X"81",X"81",X"81",X"42",X"42",X"42",X"42",X"42",X"42",X"42",X"FF",X"FF",X"FF",X"FF",X"42",X"42",
		X"00",X"00",X"00",X"0F",X"09",X"19",X"11",X"33",X"22",X"62",X"C6",X"84",X"0C",X"18",X"30",X"FF",
		X"FF",X"FF",X"1F",X"DF",X"DF",X"EF",X"EF",X"EF",X"F7",X"F7",X"07",X"FF",X"FF",X"EF",X"EF",X"EF",
		X"88",X"88",X"88",X"44",X"44",X"24",X"24",X"24",X"24",X"24",X"FF",X"FF",X"FF",X"FF",X"24",X"24",
		X"00",X"00",X"00",X"01",X"01",X"03",X"06",X"0F",X"FF",X"FF",X"F0",X"77",X"77",X"7B",X"3B",X"3D",
		X"1D",X"1E",X"0E",X"0F",X"07",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F8",X"FC",X"FE",X"FF",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"FF",X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"7F",X"3F",X"1F",X"0F",X"07",X"03",X"01",
		X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"80",
		X"C0",X"E0",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"00",X"80",X"C0",X"E0",X"F8",X"FC",X"FF",X"FF",
		X"01",X"1F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"03",X"07",X"0F",X"1F",
		X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"07",
		X"07",X"0F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"8F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"07",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"01",X"07",X"0F",X"3F",X"7F",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"F8",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"F0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"F0",X"C0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FC",X"F0",X"E0",X"E0",X"C0",X"C0",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",
		X"F8",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",
		X"F0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F0",
		X"F0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"3F",X"1F",X"1F",X"0F",X"03",X"01",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"07",X"03",X"FF",X"FF",X"E7",X"81",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"3C",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",X"1F",X"07",X"03",X"03",X"01",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FC",X"F8",X"F0",X"E0",X"C0",X"C0",X"80",X"80",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"F0",X"E0",X"C0",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7C",X"30",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"1F",X"0F",X"0F",X"07",X"07",X"03",X"03",X"01",X"01",X"00",
		X"FF",X"FF",X"FF",X"FE",X"F8",X"E0",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FE",X"FE",X"FC",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"7F",X"3F",X"1F",X"0F",X"06",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"03",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"3F",X"3F",X"3F",X"1F",X"1F",X"0F",X"07",X"03",X"01",
		X"FF",X"7F",X"7F",X"7F",X"3F",X"1F",X"1F",X"0F",X"0F",X"07",X"03",X"01",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"E1",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FC",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FC",X"F8",X"F8",X"F0",X"E0",X"C0",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"F8",X"F0",X"F0",X"E0",X"C0",X"80",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"F8",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"2F",X"07",X"03",X"01",
		X"FF",X"FF",X"FF",X"FF",X"FE",X"FC",X"FC",X"F8",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"07",X"03",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"7F",X"3F",X"1F",
		X"1F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"07",X"07",X"03",X"01",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"1F",X"07",X"03",X"03",X"03",X"01",X"01",X"FF",X"FF",X"FE",X"FE",X"FE",X"FC",X"FC",X"FC",
		X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"B0",X"10",X"FF",X"FF",X"FF",X"07",X"03",X"03",X"01",X"00",
		X"FF",X"FF",X"FF",X"FE",X"FC",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"00",X"00",X"00",X"00",X"00",
		X"FF",X"FF",X"FF",X"FE",X"F8",X"F0",X"F0",X"E0",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",
		X"3F",X"1E",X"1C",X"08",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7F",X"3F",X"0F",X"07",X"01",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"1F",X"0F",X"0F",X"07",
		X"FF",X"FF",X"FF",X"FF",X"C0",X"80",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FC",X"FC",X"F8",X"E0",X"80",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"80",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FC",X"F8",X"F0",X"E0",X"C0",X"80",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"78",X"20",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"7F",X"3F",X"0F",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"1F",X"07",X"03",X"01",X"01",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"7F",X"3F",X"0F",X"0F",X"07",X"03",X"03",X"01",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"7F",X"1F",X"0F",X"0F",X"07",X"03",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"3F",X"0F",X"00",X"00",X"FF",X"7F",X"7F",X"7F",X"3F",X"0C",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FC",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"E0",X"F0",X"F8",X"FE",X"FF",X"FF",X"FF",X"C0",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"C0",X"F0",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",
		X"F0",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"80",X"C0",
		X"C0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"80",X"80",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"E0",
		X"F0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"C0",X"E0",X"F0",X"F0",X"F0",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"E1",X"F1",X"F3",X"F3",X"FF",X"FF",X"FF",X"FF",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"6F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"03",
		X"07",X"0F",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"01",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"01",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"3F",
		X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",
		X"07",X"0F",X"0F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"81",X"C3",X"E7",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"E0",
		X"F0",X"F0",X"F8",X"FC",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"C0",X"E0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"C0",X"F0",X"F8",X"F8",X"FC",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"06",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",
		X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"FF",X"00",X"00",X"00",X"00",X"00",X"80",X"C0",X"C0",
		X"C0",X"C0",X"E0",X"F0",X"F0",X"F8",X"FE",X"FF",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"C0",X"C0",
		X"C0",X"E0",X"F0",X"F8",X"FE",X"FE",X"FC",X"FC",X"FC",X"F8",X"FC",X"FE",X"FE",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"FC",X"FE",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"80",X"E0",X"F0",X"F8",X"F8",
		X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"07",X"1F",X"7F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",
		X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"3F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",
		X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"1F",
		X"1F",X"1F",X"3F",X"3F",X"7F",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"03",X"07",X"07",X"0F",X"1F",X"3F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"03",X"07",X"0F",X"0F",X"1F",X"3F",X"7F",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"01",
		X"03",X"07",X"0F",X"3F",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"01",X"03",X"1F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FE",X"FC",X"F8",X"F8",X"F0",X"F0",X"F0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FC",X"FC",X"FC",X"FC",X"FC",
		X"FC",X"F8",X"F8",X"F8",X"F8",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"C0",X"C0",X"C0",X"80",X"80",
		X"80",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FE",X"FE",X"FE",
		X"FC",X"FC",X"FC",X"FC",X"F8",X"F8",X"F8",X"F0",X"F0",X"F0",X"F0",X"E0",X"E0",X"E0",X"E0",X"E0",
		X"C0",X"C0",X"C0",X"C0",X"80",X"80",X"00",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"7E",X"7E",X"7E",X"3E",X"3C",X"3C",X"18",X"FF",X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",
		X"3F",X"3F",X"3F",X"3F",X"1F",X"1F",X"1F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"07",X"03",X"03",
		X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"00",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"7F",X"7F",X"7F",X"3F",X"3F",X"1F",X"1F",X"1F",X"1F",X"0F",X"0F",X"07",X"07",
		X"03",X"03",X"03",X"01",X"01",X"01",X"01",X"01",X"01",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"7F",X"3F",X"3F",X"1F",X"1F",X"0F",X"0F",X"0F",X"0F",X"07",X"07",X"07",X"03",X"03",X"01",X"01",
		X"80",X"C0",X"C0",X"E0",X"F0",X"F8",X"F8",X"FE",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"80",X"C0",X"C0",X"E0",X"E0",X"F0",X"F0",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"C0",X"C0",X"C0",X"E0",X"E0",
		X"E0",X"F0",X"F0",X"F8",X"F8",X"FC",X"FC",X"FC",X"FC",X"FE",X"FE",X"FE",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"80",X"80",X"80",X"C0",X"C0",X"E0",
		X"E0",X"E0",X"F0",X"F0",X"F0",X"F8",X"F8",X"F8",X"FC",X"FC",X"FE",X"FE",X"FE",X"FE",X"FE",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"78",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"03",X"07",X"0F",X"0F",X"1F",X"1F",X"3F",X"3F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"07",X"0F",X"0F",
		X"0F",X"1F",X"1F",X"3F",X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"00",X"00",X"00",X"00",X"00",X"01",X"01",X"01",X"03",X"03",X"07",X"07",X"0F",X"0F",X"1F",X"3F",
		X"3F",X"3F",X"7F",X"7F",X"7F",X"7F",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"01",X"01",X"01",X"03",X"03",X"03",X"07",X"07",X"0F",X"0F",X"0F",X"1F",X"3F",X"7F",X"7F",X"7F",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
