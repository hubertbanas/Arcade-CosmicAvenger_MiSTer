library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu1 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu1 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"31",X"00",X"6C",X"C3",X"1E",X"01",X"FF",X"FF",X"5E",X"23",X"56",X"23",X"EB",X"C9",X"FF",X"FF",
		X"77",X"23",X"10",X"FC",X"0D",X"20",X"F9",X"C9",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"21",X"01",X"90",X"C3",X"71",X"05",X"FF",X"FF",X"F5",X"C5",X"D5",X"E5",X"C3",X"7C",X"00",X"C1",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"F5",X"C5",X"D5",X"E5",X"3A",X"03",X"90",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"CD",X"8F",X"00",X"E1",X"D1",X"C1",X"F1",X"ED",X"45",X"3A",X"03",X"90",X"E6",
		X"0F",X"C6",X"10",X"CD",X"8F",X"00",X"3A",X"00",X"80",X"E1",X"D1",X"C1",X"F1",X"FB",X"C9",X"47",
		X"3A",X"02",X"60",X"A7",X"C0",X"1E",X"06",X"CD",X"00",X"07",X"78",X"87",X"5F",X"16",X"00",X"21",
		X"DE",X"00",X"19",X"EB",X"68",X"01",X"05",X"60",X"09",X"34",X"1A",X"BE",X"C0",X"47",X"3A",X"04",
		X"60",X"4F",X"13",X"1A",X"81",X"27",X"38",X"0B",X"FE",X"99",X"28",X"07",X"32",X"04",X"60",X"36",
		X"00",X"18",X"07",X"3E",X"99",X"32",X"04",X"60",X"05",X"70",X"3A",X"00",X"60",X"17",X"D8",X"AF",
		X"32",X"45",X"63",X"32",X"46",X"63",X"21",X"47",X"63",X"CB",X"FE",X"CB",X"E6",X"C9",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"01",X"03",X"02",X"03",X"01",
		X"02",X"03",X"02",X"01",X"01",X"05",X"01",X"04",X"01",X"03",X"01",X"02",X"01",X"01",X"01",X"01",
		X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"01",X"04",X"01",X"03",X"02",X"03",X"01",
		X"02",X"03",X"02",X"01",X"01",X"05",X"01",X"04",X"01",X"03",X"01",X"02",X"01",X"01",X"3A",X"00",
		X"90",X"47",X"3A",X"01",X"90",X"A0",X"E6",X"10",X"CA",X"09",X"02",X"21",X"00",X"60",X"11",X"01",
		X"60",X"01",X"FF",X"0F",X"36",X"00",X"ED",X"B0",X"3A",X"02",X"90",X"E6",X"30",X"0F",X"0F",X"0F",
		X"47",X"0F",X"80",X"4F",X"06",X"00",X"21",X"E3",X"01",X"09",X"11",X"73",X"60",X"01",X"03",X"00",
		X"ED",X"B0",X"11",X"25",X"60",X"3E",X"05",X"21",X"73",X"60",X"01",X"03",X"00",X"ED",X"B0",X"21",
		X"FF",X"01",X"01",X"0A",X"00",X"ED",X"B0",X"3D",X"20",X"ED",X"21",X"5B",X"36",X"22",X"76",X"60",
		X"21",X"00",X"04",X"22",X"78",X"60",X"21",X"00",X"03",X"22",X"7A",X"60",X"CD",X"91",X"52",X"3A",
		X"02",X"90",X"2F",X"E6",X"03",X"32",X"DC",X"60",X"47",X"87",X"87",X"5F",X"16",X"00",X"DD",X"21",
		X"EF",X"01",X"DD",X"19",X"DD",X"6E",X"00",X"DD",X"66",X"01",X"22",X"DD",X"60",X"DD",X"6E",X"02",
		X"DD",X"66",X"03",X"22",X"DF",X"60",X"A7",X"3E",X"1E",X"28",X"02",X"3E",X"0F",X"32",X"E1",X"60",
		X"78",X"2F",X"E6",X"03",X"3E",X"3C",X"20",X"02",X"3E",X"1E",X"32",X"E2",X"60",X"78",X"21",X"00",
		X"02",X"A7",X"28",X"03",X"21",X"80",X"02",X"22",X"E3",X"60",X"21",X"00",X"01",X"E6",X"02",X"28",
		X"01",X"29",X"22",X"E5",X"60",X"3E",X"80",X"32",X"45",X"63",X"ED",X"56",X"3A",X"00",X"80",X"FB",
		X"C3",X"11",X"04",X"00",X"00",X"00",X"01",X"00",X"00",X"00",X"80",X"00",X"00",X"50",X"00",X"B4",
		X"00",X"30",X"0D",X"B4",X"00",X"30",X"0D",X"00",X"01",X"00",X"0C",X"80",X"01",X"00",X"0A",X"1E",
		X"17",X"12",X"1F",X"0E",X"1B",X"1C",X"0A",X"15",X"28",X"21",X"00",X"B0",X"36",X"9F",X"36",X"BF",
		X"36",X"DF",X"36",X"FF",X"21",X"00",X"C0",X"36",X"9F",X"36",X"BF",X"36",X"DF",X"36",X"FF",X"21",
		X"00",X"D0",X"36",X"24",X"23",X"7C",X"FE",X"E0",X"38",X"F8",X"0E",X"40",X"11",X"20",X"00",X"21",
		X"00",X"70",X"06",X"20",X"36",X"00",X"19",X"10",X"FB",X"0D",X"20",X"F3",X"DD",X"21",X"ED",X"D1",
		X"DD",X"36",X"00",X"1B",X"DD",X"36",X"01",X"18",X"DD",X"36",X"02",X"16",X"21",X"00",X"00",X"11",
		X"00",X"00",X"AF",X"06",X"10",X"86",X"2C",X"20",X"FC",X"24",X"10",X"F9",X"BB",X"28",X"10",X"16",
		X"FF",X"7B",X"C6",X"01",X"DD",X"77",X"04",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"1C",
		X"7B",X"FE",X"06",X"38",X"DD",X"CB",X"7A",X"C2",X"00",X"00",X"DD",X"36",X"04",X"18",X"DD",X"36",
		X"05",X"14",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"DD",X"36",X"00",X"1B",X"DD",X"36",
		X"01",X"0A",X"DD",X"36",X"02",X"16",X"DD",X"36",X"04",X"24",X"DD",X"36",X"05",X"24",X"1E",X"FF",
		X"21",X"00",X"60",X"16",X"10",X"7B",X"0E",X"10",X"06",X"10",X"C6",X"2F",X"77",X"23",X"10",X"FA",
		X"3D",X"0D",X"20",X"F4",X"3D",X"15",X"20",X"EE",X"21",X"00",X"60",X"16",X"10",X"7B",X"0E",X"10",
		X"06",X"10",X"C6",X"2F",X"BE",X"20",X"23",X"23",X"10",X"F8",X"3D",X"0D",X"20",X"F2",X"3D",X"15",
		X"20",X"EC",X"7B",X"D6",X"0F",X"5F",X"30",X"C8",X"DD",X"36",X"04",X"18",X"DD",X"36",X"05",X"14",
		X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"18",X"15",X"7C",X"E6",X"0C",X"0F",X"0F",X"C6",
		X"01",X"DD",X"77",X"04",X"01",X"00",X"00",X"0B",X"78",X"B1",X"20",X"FB",X"C3",X"00",X"00",X"21",
		X"34",X"03",X"CD",X"75",X"09",X"21",X"00",X"60",X"36",X"00",X"11",X"01",X"60",X"01",X"FF",X"0F",
		X"ED",X"B0",X"1E",X"00",X"D5",X"CD",X"00",X"07",X"06",X"00",X"C5",X"F7",X"CD",X"8B",X"50",X"C1",
		X"10",X"F8",X"D1",X"D5",X"CD",X"0E",X"07",X"F7",X"CD",X"8B",X"50",X"D1",X"1C",X"7B",X"FE",X"1A",
		X"38",X"E2",X"18",X"09",X"ED",X"D1",X"06",X"1C",X"18",X"1E",X"17",X"0D",X"24",X"1E",X"FF",X"21",
		X"00",X"D0",X"16",X"04",X"7B",X"0E",X"10",X"06",X"10",X"C6",X"2F",X"77",X"23",X"10",X"FA",X"3D",
		X"0D",X"20",X"F4",X"3D",X"15",X"20",X"EE",X"21",X"00",X"D0",X"16",X"04",X"7B",X"0E",X"10",X"06",
		X"10",X"C6",X"2F",X"BE",X"20",X"5F",X"23",X"10",X"F8",X"3D",X"0D",X"20",X"F2",X"3D",X"15",X"20",
		X"EC",X"7B",X"D6",X"0F",X"5F",X"30",X"C8",X"1E",X"10",X"21",X"00",X"D4",X"16",X"04",X"7B",X"0E",
		X"10",X"06",X"10",X"3C",X"77",X"23",X"10",X"FB",X"3C",X"0D",X"20",X"F5",X"3C",X"15",X"20",X"EF",
		X"21",X"00",X"D4",X"16",X"04",X"7B",X"0E",X"10",X"06",X"10",X"C5",X"3C",X"E6",X"0F",X"47",X"7E",
		X"E6",X"0F",X"B8",X"C1",X"20",X"23",X"23",X"10",X"F1",X"3C",X"0D",X"20",X"EB",X"3C",X"15",X"20",
		X"E5",X"1D",X"20",X"C5",X"AF",X"CD",X"D5",X"07",X"21",X"E0",X"03",X"CD",X"75",X"09",X"06",X"3C",
		X"F7",X"10",X"FD",X"18",X"2C",X"16",X"01",X"18",X"02",X"16",X"02",X"21",X"80",X"D0",X"01",X"00",
		X"03",X"72",X"23",X"0B",X"78",X"B1",X"20",X"F9",X"06",X"3C",X"F7",X"10",X"FD",X"C3",X"00",X"00",
		X"E9",X"D1",X"0E",X"0D",X"12",X"1C",X"19",X"15",X"0A",X"22",X"24",X"1B",X"0A",X"16",X"24",X"18",
		X"14",X"AF",X"CD",X"D5",X"07",X"21",X"03",X"04",X"CD",X"75",X"09",X"06",X"78",X"F7",X"10",X"FD",
		X"C3",X"00",X"00",X"EA",X"D1",X"0B",X"1F",X"0E",X"1B",X"1C",X"12",X"18",X"17",X"24",X"05",X"25",
		X"00",X"F7",X"FD",X"21",X"00",X"60",X"FD",X"CB",X"01",X"7E",X"C4",X"B4",X"05",X"FD",X"CB",X"01",
		X"76",X"C4",X"89",X"05",X"FD",X"CB",X"01",X"6E",X"C4",X"D8",X"06",X"FD",X"36",X"01",X"00",X"CD",
		X"8B",X"50",X"21",X"AD",X"04",X"3A",X"00",X"60",X"FD",X"21",X"E7",X"60",X"CB",X"5F",X"28",X"04",
		X"FD",X"21",X"16",X"62",X"5E",X"23",X"56",X"23",X"D5",X"DD",X"E1",X"5E",X"23",X"56",X"23",X"DD",
		X"CB",X"00",X"7E",X"28",X"17",X"DD",X"7E",X"01",X"A7",X"28",X"05",X"DD",X"35",X"01",X"18",X"0C",
		X"FD",X"E5",X"E5",X"EB",X"01",X"69",X"04",X"C5",X"E9",X"E1",X"FD",X"E1",X"EB",X"21",X"01",X"60",
		X"3A",X"01",X"90",X"07",X"2F",X"AE",X"E6",X"01",X"28",X"14",X"34",X"7E",X"E6",X"1F",X"FE",X"02",
		X"20",X"0C",X"FD",X"E5",X"D5",X"CD",X"8B",X"50",X"CD",X"79",X"05",X"D1",X"FD",X"E1",X"21",X"71",
		X"05",X"A7",X"ED",X"52",X"28",X"03",X"EB",X"18",X"AB",X"3A",X"01",X"60",X"E6",X"1F",X"FE",X"02",
		X"30",X"04",X"F7",X"CD",X"8B",X"50",X"21",X"03",X"60",X"34",X"C3",X"11",X"04",X"68",X"63",X"38",
		X"2A",X"79",X"63",X"38",X"2A",X"60",X"63",X"B8",X"29",X"54",X"63",X"59",X"26",X"8A",X"63",X"69",
		X"12",X"1C",X"65",X"4C",X"46",X"29",X"65",X"4C",X"46",X"36",X"65",X"4C",X"46",X"43",X"65",X"4C",
		X"46",X"50",X"65",X"4C",X"46",X"5D",X"65",X"4C",X"46",X"6A",X"65",X"4C",X"46",X"77",X"65",X"4C",
		X"46",X"80",X"64",X"08",X"3B",X"8A",X"64",X"08",X"3B",X"94",X"64",X"08",X"3B",X"9E",X"64",X"08",
		X"3B",X"A8",X"64",X"08",X"3B",X"B2",X"64",X"08",X"3B",X"BC",X"64",X"08",X"3B",X"C6",X"64",X"08",
		X"3B",X"FC",X"63",X"D7",X"36",X"07",X"64",X"D7",X"36",X"12",X"64",X"D7",X"36",X"1D",X"64",X"D7",
		X"36",X"28",X"64",X"D7",X"36",X"33",X"64",X"D7",X"36",X"3E",X"64",X"D7",X"36",X"49",X"64",X"D7",
		X"36",X"54",X"64",X"D7",X"36",X"5F",X"64",X"D7",X"36",X"6A",X"64",X"D7",X"36",X"75",X"64",X"D7",
		X"36",X"D0",X"64",X"96",X"40",X"DC",X"64",X"94",X"43",X"E4",X"64",X"94",X"43",X"EC",X"64",X"94",
		X"43",X"F4",X"64",X"94",X"43",X"FC",X"64",X"94",X"43",X"04",X"65",X"94",X"43",X"0C",X"65",X"94",
		X"43",X"14",X"65",X"94",X"43",X"F9",X"63",X"9A",X"35",X"EE",X"63",X"03",X"2D",X"84",X"65",X"00",
		X"2C",X"86",X"65",X"2C",X"2C",X"45",X"63",X"C4",X"0C",X"47",X"63",X"65",X"0D",X"49",X"63",X"BE",
		X"0E",X"CB",X"7E",X"20",X"FC",X"CB",X"7E",X"28",X"FC",X"21",X"02",X"60",X"7E",X"A7",X"28",X"01",
		X"35",X"3A",X"00",X"90",X"17",X"D8",X"36",X"0A",X"C9",X"21",X"00",X"71",X"0E",X"C0",X"16",X"02",
		X"1E",X"60",X"CD",X"9C",X"05",X"21",X"40",X"71",X"16",X"0B",X"1E",X"60",X"06",X"04",X"36",X"C8",
		X"23",X"71",X"23",X"72",X"23",X"73",X"23",X"79",X"C6",X"04",X"4F",X"7B",X"C6",X"10",X"5F",X"10",
		X"ED",X"36",X"00",X"C9",X"21",X"89",X"65",X"11",X"80",X"70",X"DD",X"21",X"89",X"68",X"06",X"0C",
		X"C5",X"E5",X"DD",X"7E",X"00",X"87",X"28",X"26",X"D5",X"87",X"4F",X"06",X"00",X"ED",X"B0",X"DD",
		X"36",X"00",X"00",X"FE",X"40",X"28",X"13",X"FE",X"20",X"30",X"0A",X"AF",X"12",X"D1",X"21",X"20",
		X"00",X"19",X"77",X"18",X"0F",X"AF",X"12",X"D1",X"18",X"0A",X"C1",X"C1",X"18",X"0E",X"12",X"21",
		X"20",X"00",X"19",X"77",X"E1",X"01",X"40",X"00",X"09",X"EB",X"09",X"EB",X"C1",X"DD",X"23",X"10",
		X"BF",X"C9",X"DD",X"66",X"03",X"DD",X"6E",X"05",X"3A",X"00",X"60",X"1F",X"30",X"0C",X"78",X"EE",
		X"30",X"47",X"7C",X"2F",X"3D",X"67",X"7D",X"2F",X"3D",X"6F",X"CB",X"70",X"20",X"09",X"7C",X"D6",
		X"02",X"5F",X"7D",X"D6",X"0B",X"18",X"07",X"7C",X"D6",X"06",X"5F",X"7D",X"D6",X"07",X"FE",X"D8",
		X"D0",X"D6",X"18",X"D8",X"6F",X"E6",X"0F",X"B0",X"47",X"DD",X"E5",X"D5",X"7D",X"E6",X"F0",X"6F",
		X"26",X"00",X"29",X"29",X"EB",X"DD",X"21",X"89",X"65",X"DD",X"19",X"0F",X"0F",X"0F",X"0F",X"5F",
		X"16",X"00",X"21",X"89",X"68",X"19",X"7E",X"FE",X"10",X"30",X"1B",X"87",X"87",X"5F",X"DD",X"19",
		X"D1",X"DD",X"70",X"00",X"DD",X"71",X"01",X"DD",X"72",X"02",X"DD",X"73",X"03",X"34",X"DD",X"E1",
		X"21",X"01",X"60",X"CB",X"FE",X"C9",X"D1",X"DD",X"E1",X"C9",X"DD",X"56",X"02",X"DD",X"5E",X"03",
		X"2A",X"78",X"60",X"3A",X"7B",X"60",X"AC",X"E6",X"80",X"28",X"13",X"7A",X"AC",X"E6",X"80",X"20",
		X"05",X"ED",X"52",X"30",X"12",X"C9",X"2A",X"7A",X"60",X"ED",X"52",X"38",X"0A",X"C9",X"ED",X"52",
		X"D8",X"2A",X"7A",X"60",X"ED",X"52",X"D0",X"7B",X"CB",X"1A",X"1F",X"CB",X"1A",X"1F",X"CB",X"1A",
		X"1F",X"CB",X"1A",X"1F",X"C6",X"70",X"67",X"DD",X"7E",X"05",X"D6",X"48",X"30",X"03",X"AF",X"18",
		X"0B",X"E6",X"F8",X"1F",X"1F",X"1F",X"FE",X"0E",X"38",X"02",X"3E",X"0D",X"C6",X"28",X"6F",X"50",
		X"06",X"80",X"0E",X"6E",X"CD",X"08",X"06",X"C9",X"21",X"61",X"D0",X"11",X"7F",X"60",X"FD",X"46",
		X"00",X"0E",X"12",X"1A",X"CB",X"40",X"28",X"02",X"2F",X"3D",X"77",X"0D",X"C8",X"13",X"13",X"7D",
		X"C6",X"20",X"FE",X"80",X"38",X"02",X"D6",X"7F",X"6F",X"18",X"E8",X"3A",X"00",X"60",X"17",X"D0",
		X"16",X"00",X"21",X"06",X"6C",X"19",X"36",X"01",X"21",X"C2",X"60",X"19",X"34",X"C9",X"16",X"00",
		X"21",X"C2",X"60",X"19",X"7E",X"A7",X"28",X"02",X"35",X"C0",X"21",X"06",X"6C",X"19",X"CB",X"D6",
		X"C9",X"3A",X"00",X"60",X"17",X"D0",X"FD",X"E5",X"E1",X"23",X"23",X"23",X"06",X"03",X"AF",X"1A",
		X"8E",X"27",X"77",X"1B",X"2B",X"10",X"F8",X"E5",X"CD",X"16",X"09",X"D1",X"3A",X"02",X"90",X"E6",
		X"30",X"C8",X"3E",X"04",X"21",X"00",X"60",X"CB",X"5E",X"28",X"01",X"0F",X"4F",X"A6",X"C0",X"E5",
		X"13",X"21",X"73",X"60",X"CD",X"6B",X"07",X"E1",X"D8",X"79",X"B6",X"77",X"FD",X"7E",X"00",X"FD",
		X"34",X"00",X"CD",X"AF",X"09",X"1E",X"06",X"CD",X"FB",X"06",X"C9",X"06",X"03",X"1A",X"BE",X"C0",
		X"13",X"23",X"10",X"F9",X"C9",X"2A",X"76",X"60",X"54",X"5D",X"29",X"19",X"7B",X"84",X"67",X"22",
		X"76",X"60",X"C9",X"CD",X"D5",X"07",X"21",X"89",X"68",X"11",X"8A",X"68",X"01",X"0B",X"00",X"36",
		X"00",X"ED",X"B0",X"F7",X"21",X"00",X"70",X"11",X"20",X"00",X"06",X"20",X"36",X"00",X"19",X"10",
		X"FB",X"21",X"C3",X"07",X"CD",X"75",X"09",X"CD",X"1D",X"09",X"21",X"CF",X"07",X"CD",X"75",X"09",
		X"CD",X"2D",X"09",X"3A",X"00",X"60",X"E6",X"10",X"C8",X"21",X"C9",X"07",X"CD",X"75",X"09",X"CD",
		X"25",X"09",X"C9",X"23",X"D3",X"03",X"01",X"1C",X"1D",X"43",X"D3",X"03",X"02",X"17",X"0D",X"33",
		X"D3",X"03",X"1D",X"18",X"19",X"87",X"4F",X"06",X"00",X"21",X"15",X"08",X"09",X"5E",X"23",X"56",
		X"21",X"00",X"D4",X"1A",X"A7",X"28",X"0C",X"4F",X"13",X"1A",X"13",X"D5",X"57",X"CD",X"0D",X"08",
		X"D1",X"18",X"F0",X"21",X"80",X"D0",X"01",X"80",X"03",X"16",X"24",X"CD",X"0D",X"08",X"21",X"00",
		X"D0",X"0E",X"80",X"16",X"00",X"CD",X"0D",X"08",X"21",X"7C",X"60",X"0E",X"46",X"72",X"23",X"0B",
		X"78",X"B1",X"20",X"F9",X"C9",X"25",X"08",X"40",X"08",X"69",X"08",X"88",X"08",X"C9",X"08",X"E2",
		X"08",X"E2",X"08",X"ED",X"08",X"FF",X"03",X"FF",X"03",X"C2",X"03",X"0A",X"01",X"56",X"06",X"06",
		X"00",X"0A",X"05",X"06",X"06",X"0A",X"01",X"06",X"00",X"0A",X"05",X"0B",X"00",X"A5",X"05",X"00",
		X"A7",X"01",X"39",X"06",X"07",X"01",X"39",X"03",X"07",X"01",X"39",X"05",X"07",X"01",X"39",X"04",
		X"07",X"01",X"F9",X"02",X"2A",X"01",X"56",X"06",X"06",X"00",X"0A",X"05",X"06",X"06",X"0A",X"01",
		X"06",X"00",X"0A",X"05",X"0B",X"00",X"A5",X"05",X"00",X"FF",X"03",X"FF",X"03",X"22",X"03",X"40",
		X"05",X"60",X"04",X"0A",X"01",X"56",X"06",X"06",X"00",X"0A",X"05",X"06",X"06",X"0A",X"01",X"06",
		X"00",X"0A",X"05",X"0B",X"00",X"A5",X"05",X"00",X"A7",X"01",X"39",X"06",X"07",X"01",X"39",X"03",
		X"07",X"01",X"39",X"05",X"07",X"01",X"39",X"04",X"07",X"01",X"39",X"02",X"20",X"06",X"20",X"01",
		X"1C",X"00",X"04",X"03",X"20",X"01",X"1C",X"00",X"04",X"03",X"20",X"01",X"1C",X"00",X"04",X"03",
		X"20",X"01",X"1C",X"05",X"04",X"04",X"20",X"01",X"06",X"00",X"0A",X"05",X"06",X"06",X"0A",X"01",
		X"06",X"00",X"0A",X"05",X"0B",X"00",X"A5",X"05",X"00",X"FF",X"05",X"FF",X"05",X"FF",X"05",X"23",
		X"05",X"06",X"00",X"0A",X"05",X"06",X"06",X"0A",X"01",X"06",X"00",X"0A",X"05",X"0B",X"00",X"A5",
		X"05",X"00",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"FF",X"01",X"04",X"01",X"00",X"87",X"05",X"10",
		X"04",X"09",X"05",X"07",X"05",X"10",X"04",X"09",X"05",X"07",X"05",X"10",X"04",X"09",X"05",X"FF",
		X"01",X"FF",X"01",X"42",X"01",X"06",X"00",X"0A",X"05",X"06",X"06",X"0A",X"01",X"06",X"00",X"0A",
		X"05",X"0B",X"00",X"A5",X"05",X"00",X"3A",X"00",X"60",X"CB",X"5F",X"20",X"08",X"11",X"27",X"D3",
		X"21",X"E8",X"60",X"18",X"0E",X"11",X"47",X"D3",X"21",X"17",X"62",X"18",X"06",X"11",X"37",X"D3",
		X"21",X"25",X"60",X"AF",X"06",X"06",X"ED",X"6F",X"20",X"05",X"F5",X"3E",X"24",X"18",X"05",X"CB",
		X"FF",X"F5",X"E6",X"0F",X"12",X"F1",X"13",X"CB",X"40",X"28",X"05",X"ED",X"6F",X"23",X"18",X"06",
		X"CB",X"50",X"20",X"02",X"CB",X"FF",X"10",X"DE",X"C9",X"5E",X"23",X"56",X"23",X"46",X"23",X"4E",
		X"23",X"C5",X"D5",X"7E",X"12",X"13",X"23",X"10",X"FA",X"D1",X"EB",X"01",X"20",X"00",X"09",X"EB",
		X"C1",X"0D",X"20",X"ED",X"C9",X"5E",X"23",X"56",X"23",X"46",X"23",X"7E",X"12",X"13",X"23",X"10",
		X"FA",X"C9",X"C5",X"E5",X"36",X"24",X"23",X"10",X"FB",X"E1",X"01",X"20",X"00",X"09",X"C1",X"0D",
		X"20",X"F0",X"C9",X"21",X"A6",X"09",X"CD",X"75",X"09",X"11",X"5C",X"D3",X"21",X"04",X"60",X"AF",
		X"06",X"02",X"CD",X"36",X"09",X"C9",X"55",X"D3",X"06",X"0C",X"1B",X"0E",X"0D",X"12",X"1D",X"21",
		X"D0",X"09",X"06",X"05",X"FD",X"7E",X"00",X"5E",X"23",X"56",X"23",X"EB",X"A7",X"28",X"08",X"3D",
		X"36",X"3B",X"23",X"36",X"3C",X"18",X"05",X"36",X"24",X"23",X"36",X"24",X"EB",X"10",X"E8",X"C9",
		X"C1",X"D0",X"C3",X"D0",X"C5",X"D0",X"A1",X"D0",X"A3",X"D0",X"21",X"E1",X"09",X"CD",X"59",X"09",
		X"C9",X"87",X"D0",X"10",X"03",X"45",X"46",X"46",X"46",X"46",X"46",X"46",X"4E",X"4E",X"46",X"46",
		X"46",X"46",X"46",X"46",X"47",X"48",X"4D",X"4D",X"4D",X"4D",X"4D",X"4D",X"4F",X"4F",X"4D",X"4D",
		X"4D",X"4D",X"4D",X"4D",X"49",X"4A",X"4B",X"4B",X"4B",X"4B",X"4B",X"4B",X"50",X"50",X"4B",X"4B",
		X"4B",X"4B",X"4B",X"4B",X"4C",X"FD",X"7E",X"00",X"CB",X"7F",X"C8",X"2F",X"CB",X"67",X"C9",X"E6",
		X"38",X"FE",X"10",X"28",X"04",X"38",X"02",X"E6",X"08",X"0F",X"0F",X"4F",X"06",X"00",X"21",X"33",
		X"0A",X"09",X"C9",X"03",X"03",X"07",X"07",X"0B",X"0B",X"78",X"86",X"47",X"23",X"79",X"86",X"4F",
		X"2B",X"DD",X"7E",X"02",X"FD",X"B6",X"02",X"C0",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"30",X"02",
		X"ED",X"44",X"B8",X"D0",X"DD",X"7E",X"05",X"FD",X"96",X"05",X"30",X"02",X"ED",X"44",X"B9",X"C9",
		X"DD",X"7E",X"05",X"E6",X"F8",X"5F",X"CD",X"F6",X"0A",X"DD",X"86",X"03",X"E6",X"F8",X"57",X"D5",
		X"CD",X"03",X"0B",X"E5",X"CD",X"15",X"0B",X"E1",X"D1",X"C0",X"DD",X"7E",X"03",X"80",X"FE",X"F8",
		X"30",X"1A",X"D9",X"86",X"D9",X"E6",X"F8",X"BA",X"28",X"12",X"D5",X"E5",X"7D",X"E6",X"E0",X"57",
		X"7D",X"3C",X"E6",X"1F",X"B2",X"6F",X"CD",X"15",X"0B",X"E1",X"D1",X"C0",X"DD",X"7E",X"03",X"90",
		X"FE",X"08",X"38",X"18",X"D9",X"86",X"D9",X"E6",X"F8",X"BA",X"28",X"10",X"D5",X"7D",X"E6",X"E0",
		X"57",X"7D",X"3D",X"E6",X"1F",X"B2",X"6F",X"CD",X"15",X"0B",X"D1",X"C0",X"DD",X"56",X"03",X"DD",
		X"7E",X"05",X"81",X"E6",X"F8",X"BB",X"28",X"15",X"D5",X"5F",X"D9",X"23",X"23",X"7E",X"2B",X"2B",
		X"D9",X"82",X"E6",X"F8",X"57",X"CD",X"03",X"0B",X"CD",X"15",X"0B",X"D1",X"C0",X"DD",X"7E",X"05",
		X"91",X"E6",X"F8",X"BB",X"C8",X"5F",X"D9",X"2B",X"2B",X"7E",X"D9",X"82",X"E6",X"F8",X"57",X"CD",
		X"03",X"0B",X"CD",X"15",X"0B",X"C9",X"0F",X"0F",X"D9",X"5F",X"16",X"00",X"21",X"71",X"60",X"19",
		X"7E",X"D9",X"C9",X"6B",X"26",X"00",X"29",X"29",X"7A",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"19",
		X"11",X"00",X"D0",X"19",X"C9",X"7E",X"11",X"00",X"04",X"19",X"CB",X"5E",X"21",X"3B",X"0B",X"28",
		X"03",X"21",X"5B",X"0B",X"5F",X"CB",X"3B",X"CB",X"3B",X"CB",X"3B",X"16",X"00",X"19",X"E6",X"07",
		X"57",X"3E",X"80",X"28",X"04",X"0F",X"15",X"20",X"FC",X"A6",X"C9",X"FF",X"C0",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"2F",X"FF",X"E5",X"DB",X"FE",X"DF",X"FD",X"BE",X"BF",
		X"6E",X"CF",X"FF",X"F7",X"83",X"7F",X"F7",X"DF",X"C0",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"DD",X"66",X"03",X"DD",X"6E",
		X"04",X"ED",X"5B",X"7C",X"60",X"A7",X"ED",X"52",X"DD",X"74",X"03",X"DD",X"75",X"04",X"D0",X"DD",
		X"35",X"02",X"C9",X"E6",X"0C",X"0F",X"5F",X"16",X"00",X"19",X"06",X"C0",X"4E",X"23",X"56",X"CD",
		X"02",X"06",X"C9",X"E0",X"0D",X"E4",X"0C",X"E8",X"05",X"E6",X"38",X"FE",X"10",X"28",X"18",X"38",
		X"02",X"E6",X"08",X"06",X"80",X"0E",X"70",X"16",X"01",X"CB",X"5F",X"28",X"06",X"06",X"C0",X"0E",
		X"34",X"16",X"01",X"CD",X"02",X"06",X"C9",X"21",X"E3",X"0B",X"06",X"04",X"C5",X"56",X"23",X"5E",
		X"23",X"4E",X"23",X"E5",X"CD",X"EF",X"0B",X"06",X"C0",X"16",X"01",X"CD",X"08",X"06",X"E1",X"C1",
		X"10",X"EA",X"C9",X"F8",X"08",X"40",X"F8",X"F8",X"38",X"08",X"F8",X"3C",X"08",X"08",X"44",X"DD",
		X"7E",X"03",X"82",X"67",X"DD",X"7E",X"05",X"83",X"6F",X"C9",X"AF",X"32",X"45",X"63",X"32",X"46",
		X"63",X"32",X"54",X"63",X"32",X"55",X"63",X"32",X"60",X"63",X"32",X"68",X"63",X"32",X"79",X"63",
		X"32",X"8A",X"63",X"21",X"94",X"63",X"11",X"05",X"00",X"06",X"12",X"CD",X"56",X"0C",X"32",X"EE",
		X"63",X"32",X"F9",X"63",X"21",X"FC",X"63",X"11",X"0B",X"00",X"06",X"0C",X"CD",X"56",X"0C",X"21",
		X"80",X"64",X"11",X"0A",X"00",X"06",X"08",X"CD",X"56",X"0C",X"32",X"D0",X"64",X"21",X"DC",X"64",
		X"11",X"08",X"00",X"06",X"08",X"CD",X"56",X"0C",X"32",X"84",X"65",X"32",X"86",X"65",X"21",X"1C",
		X"65",X"11",X"0D",X"00",X"06",X"08",X"77",X"19",X"10",X"FC",X"C9",X"3A",X"02",X"90",X"E6",X"C0",
		X"07",X"07",X"4F",X"06",X"00",X"21",X"6E",X"0C",X"09",X"7E",X"FD",X"77",X"00",X"C9",X"02",X"05",
		X"04",X"03",X"FD",X"E5",X"D1",X"13",X"62",X"6B",X"13",X"36",X"00",X"01",X"2D",X"01",X"ED",X"B0",
		X"FD",X"36",X"04",X"01",X"FD",X"36",X"05",X"FF",X"FD",X"36",X"08",X"01",X"FD",X"36",X"10",X"12",
		X"FD",X"36",X"13",X"01",X"FD",X"36",X"16",X"04",X"FD",X"36",X"1A",X"12",X"FD",X"36",X"1D",X"01",
		X"FD",X"36",X"20",X"01",X"01",X"11",X"1B",X"FD",X"70",X"25",X"FD",X"71",X"26",X"FD",X"36",X"27",
		X"01",X"FD",X"36",X"2A",X"0A",X"FD",X"70",X"2F",X"FD",X"71",X"30",X"FD",X"36",X"31",X"01",X"FD",
		X"36",X"34",X"07",X"C9",X"3A",X"1E",X"6C",X"A7",X"C0",X"DD",X"CB",X"00",X"6E",X"20",X"24",X"DD",
		X"CB",X"00",X"EE",X"AF",X"32",X"00",X"A0",X"CD",X"83",X"07",X"21",X"01",X"60",X"CB",X"F6",X"CD",
		X"93",X"09",X"21",X"44",X"0D",X"CD",X"75",X"09",X"21",X"52",X"0D",X"CD",X"75",X"09",X"DD",X"36",
		X"01",X"FF",X"C9",X"DD",X"CB",X"00",X"4E",X"20",X"1A",X"3E",X"01",X"CD",X"83",X"07",X"CD",X"93",
		X"09",X"CD",X"21",X"12",X"21",X"52",X"0D",X"CD",X"75",X"09",X"DD",X"36",X"01",X"FF",X"DD",X"CB",
		X"00",X"CE",X"C9",X"3E",X"07",X"CD",X"83",X"07",X"CD",X"93",X"09",X"FD",X"36",X"00",X"01",X"21",
		X"EB",X"60",X"36",X"00",X"11",X"EC",X"60",X"01",X"2A",X"01",X"ED",X"B0",X"CD",X"80",X"0C",X"CD",
		X"AF",X"09",X"CD",X"DA",X"09",X"21",X"8A",X"63",X"CB",X"FE",X"21",X"54",X"63",X"CB",X"FE",X"DD",
		X"36",X"00",X"00",X"C9",X"EA",X"D1",X"0B",X"12",X"17",X"1C",X"0E",X"1B",X"1D",X"24",X"0C",X"18",
		X"12",X"17",X"C8",X"D2",X"10",X"3A",X"24",X"1E",X"17",X"12",X"1F",X"0E",X"1B",X"1C",X"0A",X"15",
		X"24",X"01",X"09",X"08",X"01",X"DD",X"7E",X"00",X"E6",X"03",X"C2",X"52",X"0E",X"3A",X"1E",X"6C",
		X"A7",X"20",X"65",X"DD",X"CB",X"00",X"6E",X"20",X"47",X"DD",X"CB",X"00",X"EE",X"CD",X"FA",X"0B",
		X"32",X"49",X"63",X"32",X"00",X"A0",X"3A",X"00",X"60",X"E6",X"16",X"32",X"00",X"60",X"3E",X"02",
		X"CD",X"83",X"07",X"21",X"01",X"60",X"CB",X"F6",X"21",X"6C",X"0E",X"CD",X"75",X"09",X"21",X"73",
		X"0E",X"CD",X"75",X"09",X"21",X"94",X"0E",X"CD",X"75",X"09",X"21",X"52",X"0D",X"CD",X"75",X"09",
		X"CD",X"93",X"09",X"21",X"B3",X"0E",X"CD",X"75",X"09",X"13",X"3A",X"DC",X"60",X"C6",X"01",X"12",
		X"DD",X"CB",X"00",X"66",X"C4",X"93",X"09",X"DD",X"CB",X"00",X"A6",X"3A",X"04",X"60",X"FE",X"02",
		X"38",X"06",X"21",X"83",X"0E",X"CD",X"75",X"09",X"3A",X"04",X"60",X"FE",X"02",X"38",X"07",X"3A",
		X"00",X"90",X"E6",X"40",X"28",X"08",X"3A",X"00",X"90",X"E6",X"20",X"28",X"33",X"C9",X"DD",X"CB",
		X"00",X"CE",X"3E",X"90",X"32",X"00",X"60",X"21",X"04",X"60",X"7E",X"D6",X"02",X"27",X"77",X"FD",
		X"21",X"E7",X"60",X"CD",X"5B",X"0C",X"CD",X"72",X"0C",X"FD",X"21",X"16",X"62",X"CD",X"5B",X"0C",
		X"CD",X"72",X"0C",X"3E",X"04",X"CD",X"83",X"07",X"21",X"9D",X"0E",X"CD",X"75",X"09",X"18",X"20",
		X"DD",X"CB",X"00",X"C6",X"3E",X"80",X"32",X"00",X"60",X"21",X"04",X"60",X"7E",X"D6",X"01",X"27",
		X"77",X"FD",X"21",X"E7",X"60",X"CD",X"5B",X"0C",X"CD",X"72",X"0C",X"3E",X"04",X"CD",X"83",X"07",
		X"AF",X"32",X"00",X"A0",X"32",X"DA",X"60",X"1E",X"18",X"CD",X"0E",X"07",X"1E",X"17",X"CD",X"FB",
		X"06",X"C9",X"3E",X"07",X"CD",X"83",X"07",X"CD",X"AF",X"09",X"CD",X"DA",X"09",X"21",X"8A",X"63",
		X"CB",X"FE",X"21",X"54",X"63",X"CB",X"FE",X"DD",X"36",X"00",X"00",X"C9",X"EE",X"D1",X"04",X"19",
		X"1E",X"1C",X"11",X"29",X"D2",X"0D",X"18",X"17",X"15",X"22",X"24",X"01",X"24",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"29",X"D2",X"0E",X"01",X"24",X"18",X"1B",X"24",X"02",X"24",X"19",X"15",X"0A",
		X"22",X"0E",X"1B",X"1C",X"6D",X"D2",X"06",X"0B",X"1E",X"1D",X"1D",X"18",X"17",X"EC",X"D1",X"08",
		X"19",X"15",X"0A",X"22",X"0E",X"1B",X"24",X"01",X"EC",X"D1",X"08",X"19",X"15",X"0A",X"22",X"0E",
		X"1B",X"24",X"02",X"14",X"D3",X"08",X"0F",X"0A",X"0C",X"12",X"15",X"12",X"1D",X"22",X"DD",X"CB",
		X"00",X"56",X"C2",X"D3",X"0F",X"DD",X"CB",X"00",X"4E",X"C2",X"B9",X"0F",X"DD",X"CB",X"00",X"46",
		X"20",X"32",X"DD",X"CB",X"00",X"C6",X"01",X"10",X"0E",X"DD",X"70",X"02",X"DD",X"71",X"03",X"AF",
		X"DD",X"77",X"04",X"DD",X"77",X"05",X"DD",X"77",X"06",X"DD",X"77",X"07",X"DD",X"77",X"08",X"DD",
		X"36",X"0A",X"0A",X"3A",X"02",X"90",X"E6",X"04",X"20",X"04",X"DD",X"36",X"0A",X"03",X"21",X"00",
		X"60",X"CB",X"B6",X"C9",X"3A",X"60",X"63",X"17",X"D8",X"3A",X"68",X"63",X"17",X"D8",X"3A",X"79",
		X"63",X"17",X"D8",X"21",X"80",X"64",X"11",X"0A",X"00",X"06",X"08",X"CB",X"7E",X"C0",X"19",X"10",
		X"FA",X"21",X"DC",X"64",X"11",X"08",X"00",X"06",X"08",X"7E",X"2F",X"E6",X"88",X"C8",X"19",X"10",
		X"F8",X"21",X"1C",X"65",X"11",X"0D",X"00",X"06",X"08",X"CB",X"7E",X"C0",X"19",X"10",X"FA",X"CD",
		X"FA",X"0B",X"AF",X"32",X"CE",X"60",X"32",X"D0",X"60",X"32",X"D7",X"60",X"1E",X"0C",X"CD",X"0E",
		X"07",X"1E",X"0E",X"CD",X"0E",X"07",X"1E",X"15",X"CD",X"0E",X"07",X"21",X"00",X"60",X"CB",X"7E",
		X"28",X"4D",X"FD",X"7E",X"00",X"A7",X"28",X"0E",X"CB",X"66",X"28",X"1E",X"CD",X"ED",X"0F",X"1A",
		X"A7",X"C4",X"F7",X"0F",X"18",X"14",X"CD",X"09",X"10",X"21",X"00",X"60",X"CB",X"66",X"28",X"2F",
		X"CD",X"ED",X"0F",X"1A",X"A7",X"28",X"28",X"CD",X"F7",X"0F",X"3A",X"00",X"60",X"CB",X"67",X"28",
		X"15",X"3E",X"04",X"CD",X"83",X"07",X"21",X"9D",X"0E",X"3A",X"00",X"60",X"CB",X"5F",X"28",X"03",
		X"21",X"A8",X"0E",X"CD",X"75",X"09",X"DD",X"CB",X"00",X"CE",X"DD",X"36",X"01",X"3C",X"C9",X"DD",
		X"CB",X"00",X"D6",X"1E",X"18",X"CD",X"FB",X"06",X"C9",X"3E",X"07",X"CD",X"83",X"07",X"CD",X"AF",
		X"09",X"CD",X"DA",X"09",X"21",X"8A",X"63",X"CB",X"FE",X"21",X"54",X"63",X"CB",X"FE",X"DD",X"36",
		X"00",X"00",X"C9",X"21",X"45",X"63",X"3A",X"04",X"60",X"A7",X"28",X"03",X"21",X"47",X"63",X"CB",
		X"FE",X"21",X"00",X"60",X"7E",X"E6",X"16",X"77",X"DD",X"36",X"00",X"00",X"C9",X"11",X"16",X"62",
		X"CB",X"5E",X"C8",X"11",X"E7",X"60",X"C9",X"7E",X"EE",X"08",X"77",X"3A",X"02",X"90",X"E6",X"08",
		X"C8",X"7E",X"EE",X"01",X"77",X"32",X"00",X"A0",X"C9",X"21",X"25",X"60",X"FD",X"E5",X"D1",X"13",
		X"06",X"05",X"C5",X"D5",X"E5",X"CD",X"6B",X"07",X"30",X"0A",X"E1",X"11",X"0D",X"00",X"19",X"D1",
		X"C1",X"10",X"EF",X"C9",X"E1",X"D1",X"C1",X"3E",X"05",X"90",X"DD",X"77",X"09",X"EB",X"11",X"66",
		X"60",X"01",X"03",X"00",X"ED",X"B0",X"EB",X"36",X"24",X"54",X"5D",X"13",X"01",X"09",X"00",X"ED",
		X"B0",X"3E",X"03",X"CD",X"83",X"07",X"CD",X"21",X"12",X"21",X"16",X"12",X"CD",X"75",X"09",X"21",
		X"F7",X"D1",X"DD",X"7E",X"0A",X"FE",X"0A",X"28",X"03",X"21",X"F0",X"D1",X"36",X"25",X"21",X"22",
		X"D2",X"11",X"26",X"00",X"AF",X"0E",X"04",X"06",X"0D",X"77",X"3C",X"23",X"23",X"10",X"FA",X"19",
		X"0D",X"20",X"F4",X"21",X"3C",X"D2",X"11",X"3F",X"00",X"06",X"03",X"36",X"34",X"23",X"36",X"35",
		X"19",X"10",X"F8",X"36",X"36",X"23",X"36",X"37",X"3E",X"38",X"32",X"42",X"D2",X"1E",X"13",X"CD",
		X"FB",X"06",X"F7",X"DD",X"E5",X"CD",X"8B",X"50",X"DD",X"E1",X"DD",X"46",X"02",X"DD",X"4E",X"03",
		X"0B",X"DD",X"70",X"02",X"DD",X"71",X"03",X"78",X"B1",X"CA",X"8B",X"11",X"DD",X"7E",X"04",X"DD",
		X"BE",X"0A",X"30",X"19",X"DD",X"34",X"05",X"DD",X"7E",X"05",X"E6",X"07",X"20",X"0F",X"CD",X"E3",
		X"11",X"DD",X"CB",X"05",X"5E",X"28",X"04",X"36",X"39",X"18",X"02",X"36",X"24",X"DD",X"7E",X"06",
		X"A7",X"28",X"05",X"DD",X"35",X"06",X"18",X"67",X"CD",X"0A",X"12",X"CB",X"66",X"20",X"60",X"DD",
		X"36",X"06",X"20",X"DD",X"7E",X"07",X"FE",X"37",X"20",X"03",X"C3",X"8B",X"11",X"21",X"1D",X"12",
		X"06",X"03",X"BE",X"28",X"07",X"30",X"29",X"23",X"10",X"F8",X"18",X"24",X"DD",X"7E",X"04",X"A7",
		X"28",X"3D",X"DD",X"BE",X"0A",X"30",X"05",X"CD",X"E3",X"11",X"36",X"24",X"DD",X"35",X"04",X"CD",
		X"ED",X"11",X"36",X"24",X"CD",X"DE",X"11",X"36",X"24",X"1E",X"0D",X"CD",X"FB",X"06",X"18",X"1F",
		X"90",X"47",X"DD",X"7E",X"04",X"DD",X"BE",X"0A",X"30",X"15",X"CD",X"ED",X"11",X"70",X"CD",X"DE",
		X"11",X"70",X"CD",X"E3",X"11",X"36",X"24",X"DD",X"34",X"04",X"1E",X"04",X"CD",X"FB",X"06",X"DD",
		X"7E",X"08",X"A7",X"28",X"06",X"DD",X"35",X"08",X"C3",X"92",X"10",X"CD",X"0A",X"12",X"7E",X"2F",
		X"E6",X"05",X"CA",X"92",X"10",X"DD",X"36",X"08",X"06",X"CB",X"57",X"20",X"11",X"DD",X"7E",X"07",
		X"A7",X"CA",X"92",X"10",X"CD",X"F2",X"11",X"36",X"24",X"DD",X"35",X"07",X"18",X"10",X"DD",X"7E",
		X"07",X"FE",X"37",X"CA",X"92",X"10",X"CD",X"F2",X"11",X"36",X"24",X"DD",X"34",X"07",X"CD",X"F2",
		X"11",X"36",X"38",X"1E",X"0F",X"CD",X"FB",X"06",X"C3",X"92",X"10",X"DD",X"7E",X"09",X"FE",X"04",
		X"28",X"11",X"2F",X"C6",X"05",X"21",X"58",X"60",X"11",X"65",X"60",X"01",X"0D",X"00",X"ED",X"B8",
		X"3D",X"20",X"F8",X"DD",X"7E",X"09",X"4F",X"87",X"87",X"47",X"87",X"80",X"81",X"5F",X"16",X"00",
		X"21",X"25",X"60",X"19",X"EB",X"21",X"66",X"60",X"01",X"0D",X"00",X"ED",X"B0",X"3E",X"01",X"CD",
		X"83",X"07",X"CD",X"21",X"12",X"1E",X"13",X"CD",X"0E",X"07",X"1E",X"19",X"CD",X"FB",X"06",X"06",
		X"FF",X"F7",X"DD",X"E5",X"C5",X"CD",X"8B",X"50",X"C1",X"DD",X"E1",X"10",X"F4",X"C9",X"21",X"ED",
		X"D1",X"18",X"03",X"21",X"0D",X"D2",X"DD",X"5E",X"04",X"16",X"00",X"19",X"C9",X"21",X"69",X"60",
		X"18",X"F4",X"21",X"42",X"D2",X"11",X"40",X"00",X"DD",X"7E",X"07",X"06",X"03",X"FE",X"0E",X"38",
		X"05",X"D6",X"0E",X"19",X"10",X"F7",X"87",X"5F",X"19",X"C9",X"21",X"00",X"90",X"3A",X"00",X"60",
		X"1F",X"D0",X"21",X"01",X"90",X"C9",X"E8",X"D1",X"04",X"17",X"0A",X"16",X"0E",X"29",X"1B",X"0D",
		X"C9",X"21",X"4A",X"12",X"0E",X"05",X"CD",X"75",X"09",X"0D",X"20",X"FA",X"21",X"25",X"60",X"11",
		X"AA",X"D0",X"06",X"05",X"C5",X"D5",X"CD",X"33",X"09",X"13",X"06",X"0A",X"CD",X"7B",X"09",X"D1",
		X"EB",X"01",X"40",X"00",X"09",X"EB",X"C1",X"10",X"EB",X"C9",X"A5",X"D0",X"04",X"17",X"18",X"01",
		X"28",X"E5",X"D0",X"03",X"17",X"18",X"02",X"25",X"D1",X"03",X"17",X"18",X"03",X"65",X"D1",X"03",
		X"17",X"18",X"04",X"A5",X"D1",X"03",X"17",X"18",X"05",X"21",X"00",X"60",X"CB",X"76",X"C2",X"3B",
		X"13",X"21",X"54",X"63",X"CB",X"7E",X"20",X"29",X"FD",X"7E",X"0C",X"E6",X"F8",X"FD",X"77",X"0C",
		X"FD",X"36",X"0D",X"00",X"11",X"17",X"00",X"CD",X"25",X"13",X"11",X"21",X"00",X"CD",X"25",X"13",
		X"11",X"2B",X"00",X"CD",X"25",X"13",X"11",X"35",X"00",X"CD",X"25",X"13",X"DD",X"36",X"00",X"00",
		X"C9",X"DD",X"CB",X"00",X"6E",X"20",X"4C",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"02",X"00",X"DD",
		X"36",X"03",X"00",X"DD",X"36",X"09",X"00",X"21",X"00",X"04",X"22",X"7C",X"60",X"21",X"7E",X"60",
		X"36",X"00",X"11",X"7F",X"60",X"01",X"23",X"00",X"ED",X"B0",X"DD",X"E5",X"DD",X"21",X"94",X"63",
		X"11",X"05",X"00",X"06",X"12",X"DD",X"36",X"00",X"00",X"DD",X"36",X"03",X"00",X"DD",X"19",X"10",
		X"F4",X"DD",X"E1",X"21",X"EE",X"63",X"CB",X"FE",X"21",X"F9",X"63",X"CB",X"FE",X"21",X"84",X"65",
		X"CB",X"FE",X"C9",X"3A",X"A1",X"60",X"DD",X"96",X"09",X"FE",X"08",X"38",X"12",X"CD",X"0B",X"14",
		X"CD",X"A9",X"18",X"3A",X"A1",X"60",X"DD",X"77",X"09",X"CD",X"81",X"19",X"CD",X"81",X"19",X"21",
		X"7F",X"60",X"06",X"12",X"7E",X"C6",X"04",X"77",X"23",X"23",X"10",X"F8",X"CD",X"C3",X"1A",X"21",
		X"01",X"60",X"CB",X"EE",X"C9",X"FD",X"E5",X"E1",X"19",X"7E",X"E6",X"F8",X"BE",X"28",X"08",X"C6",
		X"08",X"77",X"30",X"03",X"2B",X"34",X"23",X"23",X"36",X"00",X"C9",X"DD",X"CB",X"00",X"4E",X"20",
		X"1F",X"3A",X"A1",X"60",X"DD",X"96",X"09",X"FE",X"08",X"38",X"15",X"CD",X"0B",X"14",X"DD",X"CB",
		X"00",X"56",X"C4",X"30",X"18",X"CD",X"A9",X"18",X"3A",X"A1",X"60",X"E6",X"F8",X"DD",X"77",X"09",
		X"CD",X"81",X"19",X"0E",X"00",X"DD",X"7E",X"00",X"E6",X"18",X"20",X"1C",X"FD",X"7E",X"38",X"E6",
		X"60",X"20",X"15",X"21",X"A2",X"60",X"06",X"20",X"3E",X"1F",X"BE",X"38",X"05",X"7E",X"FE",X"07",
		X"28",X"03",X"23",X"10",X"F5",X"D6",X"07",X"4F",X"DD",X"E5",X"DD",X"21",X"7E",X"60",X"3E",X"00",
		X"B9",X"30",X"28",X"47",X"3E",X"12",X"90",X"87",X"87",X"87",X"5F",X"16",X"00",X"2A",X"7C",X"60",
		X"ED",X"52",X"DD",X"56",X"01",X"DD",X"5E",X"00",X"19",X"DD",X"74",X"01",X"DD",X"75",X"00",X"78",
		X"DD",X"23",X"DD",X"23",X"3C",X"FE",X"12",X"38",X"D7",X"18",X"1A",X"ED",X"5B",X"7C",X"60",X"DD",
		X"66",X"01",X"DD",X"6E",X"00",X"19",X"DD",X"74",X"01",X"DD",X"75",X"00",X"DD",X"23",X"DD",X"23",
		X"3C",X"FE",X"12",X"38",X"EA",X"DD",X"E1",X"CD",X"C3",X"1A",X"21",X"01",X"60",X"CB",X"EE",X"2A",
		X"7C",X"60",X"FD",X"56",X"0C",X"FD",X"5E",X"0D",X"19",X"FD",X"74",X"0C",X"FD",X"75",X"0D",X"D0",
		X"FD",X"66",X"0A",X"FD",X"6E",X"0B",X"23",X"FD",X"74",X"0A",X"FD",X"75",X"0B",X"FD",X"7E",X"0E",
		X"C6",X"01",X"27",X"FD",X"77",X"0E",X"FD",X"36",X"0F",X"01",X"C9",X"FD",X"CB",X"04",X"46",X"28",
		X"71",X"FD",X"CB",X"04",X"86",X"FD",X"35",X"08",X"20",X"3C",X"FD",X"34",X"05",X"FD",X"7E",X"05",
		X"FE",X"12",X"38",X"04",X"AF",X"FD",X"77",X"05",X"5F",X"16",X"00",X"21",X"F2",X"1A",X"19",X"7E",
		X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"ED",X"44",X"FD",X"77",X"09",X"7E",X"E6",X"0F",X"87",X"6F",
		X"26",X"00",X"11",X"04",X"1B",X"19",X"5E",X"23",X"56",X"1A",X"FD",X"77",X"08",X"13",X"FD",X"72",
		X"06",X"FD",X"73",X"07",X"18",X"03",X"CD",X"50",X"16",X"FD",X"E5",X"E1",X"01",X"38",X"00",X"09",
		X"CD",X"60",X"16",X"FD",X"7E",X"38",X"FE",X"A5",X"20",X"05",X"3E",X"84",X"32",X"86",X"65",X"FD",
		X"CB",X"38",X"7E",X"28",X"0D",X"CD",X"50",X"16",X"FD",X"E5",X"E1",X"01",X"4B",X"00",X"09",X"CD",
		X"60",X"16",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"11",X"38",X"00",X"DD",X"19",X"01",X"12",X"07",
		X"DD",X"CB",X"00",X"7E",X"28",X"03",X"01",X"0A",X"0F",X"DD",X"70",X"0C",X"DD",X"71",X"0D",X"DD",
		X"7E",X"00",X"E6",X"60",X"0F",X"0F",X"0F",X"F6",X"10",X"47",X"DD",X"7E",X"05",X"E6",X"E1",X"B0",
		X"47",X"CB",X"50",X"28",X"24",X"CB",X"58",X"20",X"0D",X"DD",X"7E",X"0A",X"A7",X"20",X"16",X"FD",
		X"B6",X"55",X"20",X"15",X"18",X"0B",X"FD",X"7E",X"55",X"A7",X"20",X"09",X"DD",X"B6",X"0A",X"20",
		X"08",X"3E",X"0C",X"18",X"02",X"3E",X"04",X"A8",X"47",X"DD",X"70",X"05",X"DD",X"66",X"03",X"DD",
		X"6E",X"04",X"CB",X"7E",X"28",X"53",X"7E",X"E6",X"E0",X"47",X"E6",X"60",X"20",X"0B",X"DD",X"7E",
		X"06",X"FE",X"77",X"28",X"04",X"78",X"F6",X"60",X"47",X"FD",X"70",X"5E",X"7E",X"E6",X"1F",X"FD",
		X"86",X"09",X"FD",X"77",X"5F",X"23",X"7E",X"FD",X"86",X"09",X"FD",X"77",X"60",X"23",X"E5",X"FD",
		X"7E",X"5E",X"E6",X"60",X"0F",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"9D",X"25",X"19",X"5E",
		X"23",X"56",X"1A",X"FD",X"77",X"63",X"13",X"1A",X"FD",X"77",X"64",X"13",X"FD",X"72",X"61",X"FD",
		X"73",X"62",X"E1",X"DD",X"74",X"03",X"DD",X"75",X"04",X"7E",X"47",X"E6",X"1F",X"FD",X"86",X"09",
		X"4F",X"78",X"E6",X"E0",X"B1",X"DD",X"77",X"0B",X"23",X"7E",X"DD",X"77",X"0E",X"FD",X"CB",X"5E",
		X"7E",X"28",X"03",X"FD",X"4E",X"5F",X"3A",X"A1",X"60",X"E6",X"F8",X"0F",X"0F",X"0F",X"5F",X"16",
		X"00",X"21",X"A2",X"60",X"19",X"71",X"FD",X"CB",X"5E",X"7E",X"C4",X"C0",X"17",X"CD",X"C4",X"16",
		X"DD",X"66",X"10",X"DD",X"6E",X"07",X"2B",X"DD",X"74",X"10",X"DD",X"75",X"07",X"DD",X"66",X"12",
		X"DD",X"6E",X"09",X"2B",X"DD",X"74",X"12",X"DD",X"75",X"09",X"DD",X"7E",X"0A",X"A7",X"28",X"03",
		X"DD",X"35",X"0A",X"DD",X"7E",X"07",X"DD",X"B6",X"10",X"20",X"06",X"FD",X"CB",X"04",X"C6",X"18",
		X"20",X"DD",X"7E",X"09",X"DD",X"B6",X"12",X"20",X"18",X"DD",X"7E",X"01",X"DD",X"77",X"03",X"DD",
		X"7E",X"02",X"DD",X"77",X"04",X"DD",X"7E",X"08",X"DD",X"77",X"09",X"DD",X"7E",X"11",X"DD",X"77",
		X"12",X"DD",X"E1",X"FD",X"CB",X"38",X"7E",X"C8",X"DD",X"E5",X"FD",X"E5",X"DD",X"E1",X"11",X"4B",
		X"00",X"DD",X"19",X"DD",X"36",X"0C",X"07",X"DD",X"36",X"0D",X"0B",X"DD",X"7E",X"00",X"E6",X"60",
		X"0F",X"0F",X"0F",X"47",X"DD",X"7E",X"05",X"E6",X"E1",X"B0",X"47",X"DD",X"66",X"03",X"DD",X"6E",
		X"04",X"7E",X"E6",X"1F",X"20",X"0A",X"CB",X"E0",X"23",X"DD",X"74",X"03",X"DD",X"75",X"04",X"2B",
		X"CB",X"50",X"28",X"24",X"CB",X"58",X"20",X"0D",X"FD",X"7E",X"42",X"A7",X"20",X"16",X"DD",X"B6",
		X"0A",X"20",X"15",X"18",X"0B",X"DD",X"7E",X"0A",X"A7",X"20",X"09",X"FD",X"B6",X"42",X"20",X"08",
		X"3E",X"0C",X"18",X"02",X"3E",X"04",X"A8",X"47",X"DD",X"70",X"05",X"7E",X"DD",X"77",X"0B",X"23",
		X"7E",X"DD",X"77",X"0E",X"CD",X"C4",X"16",X"DD",X"7E",X"0A",X"A7",X"28",X"03",X"DD",X"35",X"0A",
		X"DD",X"E1",X"DD",X"CB",X"00",X"E6",X"2A",X"A0",X"60",X"DD",X"74",X"04",X"DD",X"75",X"05",X"C9",
		X"FD",X"56",X"06",X"FD",X"5E",X"07",X"13",X"13",X"13",X"FD",X"72",X"06",X"FD",X"73",X"07",X"C9",
		X"1A",X"77",X"DD",X"E5",X"E5",X"DD",X"E1",X"13",X"1A",X"DD",X"77",X"05",X"13",X"1A",X"DD",X"77",
		X"06",X"DD",X"7E",X"00",X"E6",X"1F",X"87",X"4F",X"06",X"00",X"21",X"82",X"1B",X"09",X"5E",X"23",
		X"56",X"1A",X"DD",X"77",X"10",X"13",X"1A",X"DD",X"77",X"07",X"13",X"1A",X"DD",X"77",X"11",X"DD",
		X"77",X"12",X"13",X"1A",X"DD",X"77",X"08",X"DD",X"77",X"09",X"13",X"DD",X"CB",X"00",X"6E",X"28",
		X"14",X"DD",X"CB",X"00",X"76",X"20",X"08",X"1A",X"DD",X"77",X"0A",X"13",X"13",X"18",X"06",X"13",
		X"1A",X"DD",X"77",X"0A",X"13",X"DD",X"72",X"01",X"DD",X"73",X"02",X"DD",X"72",X"03",X"DD",X"73",
		X"04",X"DD",X"E1",X"C9",X"DD",X"7E",X"0B",X"E6",X"1F",X"DD",X"BE",X"0C",X"20",X"59",X"CD",X"AF",
		X"17",X"DD",X"7E",X"0B",X"E6",X"1F",X"F6",X"80",X"77",X"DD",X"7E",X"05",X"23",X"07",X"07",X"07",
		X"47",X"CD",X"86",X"17",X"70",X"23",X"DD",X"7E",X"0E",X"DD",X"86",X"06",X"77",X"DD",X"56",X"03",
		X"DD",X"5E",X"04",X"13",X"13",X"DD",X"72",X"03",X"DD",X"73",X"04",X"DD",X"CB",X"0B",X"6E",X"20",
		X"06",X"DD",X"CB",X"05",X"A6",X"18",X"04",X"DD",X"CB",X"05",X"E6",X"DD",X"CB",X"0B",X"76",X"28",
		X"6B",X"1A",X"47",X"E6",X"1F",X"FD",X"86",X"09",X"4F",X"78",X"E6",X"E0",X"B1",X"DD",X"77",X"0B",
		X"13",X"1A",X"DD",X"77",X"0E",X"18",X"55",X"DD",X"CB",X"05",X"66",X"20",X"1E",X"CD",X"AF",X"17",
		X"DD",X"7E",X"0C",X"E6",X"1F",X"F6",X"80",X"77",X"23",X"DD",X"7E",X"05",X"07",X"07",X"07",X"47",
		X"CD",X"86",X"17",X"70",X"23",X"DD",X"7E",X"06",X"77",X"18",X"31",X"CD",X"AF",X"17",X"CB",X"7E",
		X"20",X"2A",X"DD",X"7E",X"05",X"E6",X"0C",X"28",X"0B",X"FE",X"08",X"28",X"11",X"DD",X"7E",X"0C",
		X"FE",X"10",X"30",X"0A",X"DD",X"7E",X"0C",X"E6",X"1F",X"F6",X"A0",X"77",X"18",X"0E",X"DD",X"7E",
		X"0C",X"E6",X"1F",X"F6",X"80",X"77",X"23",X"36",X"06",X"23",X"36",X"FF",X"DD",X"34",X"0C",X"DD",
		X"35",X"0D",X"C2",X"C4",X"16",X"C9",X"DD",X"7E",X"00",X"E6",X"60",X"C8",X"FE",X"40",X"C8",X"78",
		X"E6",X"60",X"28",X"0D",X"FE",X"40",X"28",X"10",X"DD",X"7E",X"0B",X"E6",X"1F",X"FE",X"10",X"30",
		X"07",X"78",X"E6",X"F8",X"F6",X"07",X"47",X"C9",X"78",X"E6",X"F8",X"F6",X"06",X"47",X"C9",X"DD",
		X"7E",X"0C",X"D6",X"07",X"57",X"87",X"87",X"82",X"5F",X"16",X"00",X"21",X"94",X"63",X"19",X"C9",
		X"FD",X"66",X"61",X"FD",X"6E",X"62",X"7E",X"FD",X"77",X"65",X"E6",X"1F",X"FD",X"86",X"5F",X"FD",
		X"77",X"68",X"E5",X"F5",X"CD",X"B2",X"17",X"F1",X"F6",X"80",X"77",X"D1",X"23",X"13",X"1A",X"E6",
		X"E0",X"FD",X"B6",X"63",X"07",X"07",X"07",X"77",X"FD",X"77",X"66",X"23",X"1A",X"E6",X"1F",X"FD",
		X"86",X"64",X"77",X"FD",X"77",X"67",X"13",X"FD",X"72",X"61",X"FD",X"73",X"62",X"FD",X"7E",X"65",
		X"CB",X"7F",X"20",X"27",X"CB",X"77",X"C8",X"CB",X"6F",X"28",X"B5",X"FD",X"34",X"68",X"FD",X"7E",
		X"68",X"FD",X"BE",X"60",X"28",X"01",X"D0",X"F5",X"CD",X"B2",X"17",X"F1",X"F6",X"80",X"77",X"23",
		X"FD",X"7E",X"66",X"77",X"23",X"FD",X"7E",X"67",X"77",X"18",X"E0",X"FD",X"36",X"5E",X"00",X"C9",
		X"06",X"07",X"DD",X"7E",X"07",X"B8",X"38",X"2F",X"47",X"CD",X"B2",X"17",X"78",X"F6",X"80",X"77",
		X"23",X"36",X"02",X"23",X"36",X"40",X"04",X"11",X"03",X"00",X"19",X"3C",X"77",X"23",X"36",X"02",
		X"23",X"36",X"41",X"04",X"DD",X"35",X"07",X"DD",X"35",X"07",X"DD",X"7E",X"06",X"A7",X"20",X"07",
		X"1E",X"0C",X"CD",X"FB",X"06",X"18",X"31",X"78",X"CD",X"B2",X"17",X"78",X"DD",X"BE",X"08",X"30",
		X"10",X"F6",X"80",X"77",X"23",X"36",X"02",X"23",X"36",X"42",X"11",X"03",X"00",X"19",X"04",X"18",
		X"EA",X"F6",X"80",X"77",X"23",X"36",X"02",X"23",X"36",X"43",X"DD",X"35",X"08",X"DD",X"7E",X"08",
		X"FE",X"07",X"30",X"04",X"DD",X"CB",X"00",X"96",X"DD",X"CB",X"00",X"DE",X"2A",X"A0",X"60",X"DD",
		X"74",X"04",X"DD",X"75",X"05",X"DD",X"34",X"06",X"C9",X"2A",X"A0",X"60",X"DD",X"56",X"02",X"DD",
		X"5E",X"03",X"DD",X"74",X"02",X"DD",X"75",X"03",X"A7",X"ED",X"52",X"EB",X"DD",X"E5",X"FD",X"E5",
		X"DD",X"E1",X"01",X"10",X"00",X"DD",X"09",X"06",X"04",X"D5",X"DD",X"66",X"07",X"DD",X"6E",X"08",
		X"A7",X"ED",X"52",X"DD",X"74",X"07",X"DD",X"75",X"08",X"D2",X"74",X"19",X"DD",X"35",X"06",X"DD",
		X"CB",X"06",X"7E",X"CA",X"74",X"19",X"DD",X"CB",X"00",X"FE",X"DD",X"35",X"03",X"20",X"3F",X"DD",
		X"34",X"00",X"DD",X"7E",X"00",X"E6",X"7F",X"FE",X"12",X"38",X"05",X"DD",X"36",X"00",X"80",X"AF",
		X"5F",X"16",X"00",X"21",X"F2",X"1A",X"19",X"7E",X"E6",X"F0",X"0F",X"0F",X"0F",X"0F",X"ED",X"44",
		X"DD",X"77",X"09",X"7E",X"E6",X"0F",X"87",X"5F",X"16",X"00",X"21",X"04",X"1B",X"19",X"5E",X"23",
		X"56",X"1A",X"DD",X"77",X"03",X"13",X"DD",X"72",X"01",X"DD",X"73",X"02",X"18",X"0F",X"DD",X"56",
		X"01",X"DD",X"5E",X"02",X"13",X"13",X"13",X"DD",X"72",X"01",X"DD",X"73",X"02",X"1A",X"DD",X"77",
		X"04",X"CB",X"7F",X"28",X"0D",X"13",X"13",X"13",X"1A",X"DD",X"77",X"05",X"DD",X"72",X"01",X"DD",
		X"73",X"02",X"E6",X"1F",X"87",X"5F",X"16",X"00",X"21",X"82",X"1B",X"19",X"5E",X"23",X"56",X"EB",
		X"56",X"23",X"5E",X"EB",X"29",X"29",X"29",X"DD",X"56",X"06",X"DD",X"5E",X"07",X"19",X"DD",X"74",
		X"06",X"DD",X"75",X"07",X"11",X"0A",X"00",X"DD",X"19",X"D1",X"05",X"C2",X"C9",X"18",X"DD",X"E1",
		X"C9",X"DD",X"E5",X"DD",X"7E",X"00",X"DD",X"21",X"94",X"63",X"CB",X"47",X"28",X"04",X"DD",X"21",
		X"C1",X"63",X"06",X"09",X"C5",X"DD",X"CB",X"00",X"7E",X"C4",X"B6",X"19",X"11",X"05",X"00",X"DD",
		X"19",X"C1",X"10",X"F0",X"DD",X"E1",X"DD",X"7E",X"00",X"EE",X"01",X"DD",X"77",X"00",X"E6",X"01",
		X"C0",X"DD",X"CB",X"00",X"8E",X"C9",X"DD",X"7E",X"00",X"E6",X"1F",X"FE",X"18",X"20",X"55",X"FD",
		X"7E",X"0F",X"A7",X"28",X"4F",X"FE",X"01",X"20",X"29",X"FD",X"34",X"0F",X"FD",X"7E",X"0E",X"E6",
		X"F0",X"28",X"41",X"0F",X"0F",X"0F",X"0F",X"F5",X"CD",X"7F",X"1A",X"CD",X"8F",X"1A",X"CD",X"A6",
		X"1A",X"F1",X"77",X"7C",X"C6",X"04",X"67",X"DD",X"7E",X"01",X"E6",X"07",X"77",X"DD",X"36",X"00",
		X"00",X"C9",X"CD",X"7F",X"1A",X"CD",X"8F",X"1A",X"CD",X"A6",X"1A",X"FD",X"7E",X"0E",X"E6",X"0F",
		X"77",X"7C",X"C6",X"04",X"67",X"DD",X"7E",X"01",X"E6",X"07",X"77",X"FD",X"36",X"0F",X"00",X"DD",
		X"36",X"00",X"00",X"C9",X"DD",X"CB",X"00",X"6E",X"20",X"1A",X"CD",X"7F",X"1A",X"CD",X"8F",X"1A",
		X"CD",X"A6",X"1A",X"DD",X"7E",X"02",X"77",X"7C",X"C6",X"04",X"67",X"DD",X"7E",X"01",X"77",X"DD",
		X"36",X"00",X"00",X"C9",X"CD",X"7F",X"1A",X"7E",X"DD",X"96",X"03",X"FE",X"08",X"D8",X"7E",X"CD",
		X"A6",X"1A",X"DD",X"7E",X"04",X"A7",X"20",X"27",X"E5",X"CD",X"75",X"07",X"E1",X"E6",X"07",X"47",
		X"C6",X"51",X"77",X"7C",X"C6",X"04",X"67",X"70",X"DD",X"7E",X"00",X"E6",X"1F",X"D6",X"07",X"5F",
		X"16",X"00",X"21",X"E0",X"1A",X"19",X"7E",X"DD",X"77",X"04",X"DD",X"36",X"00",X"00",X"C9",X"DD",
		X"35",X"04",X"36",X"FF",X"7C",X"C6",X"04",X"67",X"36",X"07",X"DD",X"36",X"00",X"00",X"C9",X"DD",
		X"7E",X"00",X"E6",X"1F",X"D6",X"07",X"87",X"5F",X"16",X"00",X"21",X"7F",X"60",X"19",X"C9",X"46",
		X"3A",X"A1",X"60",X"E6",X"07",X"4F",X"78",X"E6",X"07",X"91",X"4F",X"78",X"91",X"77",X"47",X"2B",
		X"3A",X"A0",X"60",X"77",X"78",X"C9",X"E6",X"F8",X"DD",X"77",X"03",X"0F",X"0F",X"0F",X"21",X"00",
		X"D0",X"85",X"6F",X"EB",X"DD",X"7E",X"00",X"E6",X"1F",X"6F",X"26",X"00",X"29",X"29",X"29",X"29",
		X"29",X"19",X"C9",X"DD",X"7E",X"00",X"E6",X"18",X"C8",X"3A",X"A1",X"60",X"DD",X"96",X"04",X"FE",
		X"F8",X"D8",X"DD",X"7E",X"00",X"E6",X"E7",X"DD",X"77",X"00",X"1E",X"0C",X"CD",X"0E",X"07",X"C9",
		X"01",X"03",X"05",X"07",X"09",X"0B",X"0D",X"0F",X"11",X"13",X"15",X"17",X"19",X"1B",X"1D",X"1F",
		X"21",X"23",X"00",X"02",X"03",X"04",X"21",X"14",X"42",X"03",X"05",X"40",X"82",X"03",X"24",X"61",
		X"34",X"C2",X"03",X"05",X"10",X"1B",X"14",X"1B",X"18",X"1B",X"55",X"1B",X"77",X"1B",X"7B",X"1B",
		X"01",X"00",X"A0",X"77",X"01",X"00",X"20",X"AC",X"14",X"01",X"20",X"7E",X"02",X"20",X"7E",X"03",
		X"20",X"7E",X"04",X"20",X"7E",X"01",X"20",X"7E",X"02",X"20",X"7E",X"03",X"20",X"7E",X"04",X"20",
		X"7E",X"01",X"20",X"7E",X"02",X"20",X"7E",X"03",X"20",X"7E",X"04",X"20",X"7E",X"01",X"20",X"7E",
		X"02",X"20",X"7E",X"03",X"20",X"7E",X"04",X"20",X"7E",X"01",X"20",X"7E",X"02",X"20",X"7E",X"03",
		X"20",X"7E",X"04",X"20",X"7E",X"06",X"A5",X"00",X"A5",X"26",X"00",X"9B",X"C7",X"C0",X"A5",X"48",
		X"C0",X"9B",X"49",X"C0",X"A5",X"CA",X"C0",X"A5",X"4B",X"C0",X"9B",X"CC",X"C0",X"A5",X"4D",X"C0",
		X"9B",X"EE",X"00",X"A5",X"6F",X"00",X"9B",X"01",X"10",X"60",X"C6",X"01",X"91",X"20",X"E5",X"12",
		X"20",X"E5",X"A8",X"1B",X"42",X"1E",X"48",X"1E",X"52",X"1E",X"5E",X"1E",X"68",X"1E",X"A8",X"1E",
		X"F8",X"1E",X"84",X"1F",X"2E",X"20",X"A2",X"20",X"42",X"21",X"EB",X"21",X"FF",X"21",X"15",X"22",
		X"3D",X"22",X"6F",X"22",X"15",X"25",X"59",X"25",X"01",X"40",X"01",X"40",X"18",X"00",X"18",X"00",
		X"17",X"01",X"16",X"01",X"15",X"01",X"15",X"00",X"14",X"01",X"13",X"01",X"12",X"01",X"12",X"02",
		X"13",X"05",X"13",X"06",X"14",X"00",X"14",X"02",X"15",X"02",X"16",X"00",X"15",X"01",X"14",X"03",
		X"14",X"04",X"14",X"00",X"13",X"01",X"13",X"02",X"14",X"02",X"15",X"02",X"16",X"02",X"91",X"17",
		X"17",X"02",X"18",X"00",X"18",X"00",X"18",X"00",X"16",X"01",X"15",X"01",X"15",X"02",X"16",X"02",
		X"16",X"01",X"15",X"01",X"14",X"01",X"13",X"01",X"13",X"02",X"14",X"00",X"16",X"02",X"17",X"02",
		X"18",X"00",X"17",X"01",X"16",X"00",X"15",X"01",X"13",X"01",X"12",X"01",X"11",X"01",X"10",X"00",
		X"13",X"02",X"D3",X"17",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",
		X"18",X"00",X"17",X"03",X"17",X"04",X"16",X"03",X"16",X"04",X"16",X"00",X"16",X"00",X"15",X"03",
		X"15",X"04",X"14",X"03",X"14",X"04",X"14",X"00",X"14",X"00",X"13",X"03",X"13",X"04",X"12",X"03",
		X"12",X"04",X"12",X"00",X"11",X"01",X"10",X"01",X"10",X"02",X"11",X"02",X"12",X"05",X"12",X"06",
		X"13",X"00",X"13",X"02",X"14",X"02",X"91",X"17",X"15",X"02",X"18",X"00",X"18",X"00",X"18",X"00",
		X"15",X"01",X"14",X"01",X"14",X"00",X"13",X"03",X"13",X"04",X"12",X"01",X"11",X"01",X"12",X"02",
		X"13",X"02",X"14",X"02",X"15",X"02",X"90",X"17",X"16",X"02",X"18",X"00",X"18",X"00",X"18",X"00",
		X"17",X"01",X"92",X"17",X"17",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"16",X"01",X"15",X"01",
		X"14",X"01",X"13",X"01",X"13",X"02",X"14",X"00",X"14",X"05",X"14",X"06",X"15",X"05",X"15",X"06",
		X"15",X"01",X"14",X"01",X"14",X"02",X"15",X"02",X"16",X"02",X"12",X"03",X"12",X"04",X"18",X"00",
		X"12",X"03",X"12",X"04",X"17",X"00",X"13",X"05",X"13",X"06",X"18",X"00",X"14",X"05",X"14",X"06",
		X"16",X"01",X"15",X"01",X"15",X"02",X"16",X"00",X"15",X"01",X"14",X"01",X"13",X"01",X"13",X"02",
		X"14",X"02",X"15",X"02",X"16",X"02",X"17",X"00",X"17",X"00",X"90",X"17",X"17",X"02",X"18",X"00",
		X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"14",X"01",X"14",X"02",X"15",X"02",
		X"16",X"00",X"16",X"02",X"17",X"02",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",
		X"14",X"01",X"13",X"01",X"13",X"00",X"12",X"01",X"12",X"02",X"13",X"02",X"14",X"00",X"D3",X"17",
		X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"03",
		X"17",X"04",X"16",X"03",X"16",X"04",X"16",X"00",X"16",X"00",X"15",X"03",X"15",X"04",X"14",X"03",
		X"14",X"04",X"14",X"00",X"14",X"00",X"13",X"03",X"13",X"04",X"12",X"03",X"12",X"04",X"11",X"01",
		X"10",X"01",X"0F",X"01",X"10",X"01",X"15",X"02",X"91",X"17",X"16",X"02",X"18",X"00",X"18",X"00",
		X"18",X"00",X"16",X"01",X"16",X"00",X"15",X"01",X"14",X"01",X"13",X"01",X"12",X"01",X"12",X"02",
		X"13",X"02",X"14",X"02",X"15",X"00",X"15",X"02",X"16",X"00",X"16",X"05",X"16",X"06",X"17",X"05",
		X"17",X"06",X"18",X"00",X"17",X"01",X"16",X"01",X"16",X"00",X"15",X"01",X"14",X"01",X"14",X"00",
		X"13",X"01",X"12",X"01",X"12",X"02",X"13",X"02",X"14",X"02",X"91",X"15",X"15",X"02",X"16",X"00",
		X"16",X"00",X"16",X"00",X"16",X"02",X"17",X"02",X"93",X"17",X"18",X"00",X"18",X"00",X"18",X"00",
		X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"15",X"02",X"16",X"02",X"16",X"01",X"15",X"01",
		X"14",X"01",X"13",X"01",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"00",X"13",X"02",
		X"14",X"00",X"14",X"00",X"D3",X"17",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",
		X"17",X"03",X"17",X"04",X"16",X"03",X"16",X"04",X"16",X"00",X"16",X"00",X"15",X"03",X"15",X"04",
		X"14",X"03",X"14",X"04",X"14",X"00",X"14",X"00",X"13",X"03",X"13",X"04",X"12",X"03",X"12",X"04",
		X"12",X"00",X"11",X"01",X"11",X"02",X"12",X"02",X"13",X"02",X"13",X"01",X"13",X"02",X"14",X"02",
		X"16",X"01",X"16",X"00",X"16",X"02",X"17",X"02",X"17",X"01",X"16",X"01",X"15",X"01",X"12",X"01",
		X"12",X"02",X"14",X"01",X"14",X"02",X"16",X"01",X"16",X"02",X"18",X"00",X"18",X"00",X"17",X"01",
		X"16",X"01",X"13",X"03",X"13",X"04",X"13",X"02",X"15",X"01",X"15",X"02",X"16",X"02",X"17",X"00",
		X"17",X"02",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"15",X"02",X"16",X"02",
		X"17",X"02",X"00",X"1E",X"00",X"01",X"18",X"00",X"00",X"02",X"00",X"02",X"17",X"01",X"56",X"01",
		X"17",X"02",X"00",X"1E",X"00",X"02",X"56",X"03",X"17",X"04",X"56",X"05",X"17",X"06",X"00",X"02",
		X"00",X"02",X"56",X"07",X"17",X"08",X"17",X"07",X"00",X"1D",X"00",X"1D",X"0B",X"00",X"17",X"01",
		X"14",X"01",X"13",X"01",X"12",X"02",X"15",X"02",X"17",X"00",X"15",X"01",X"13",X"01",X"11",X"01",
		X"0F",X"01",X"0F",X"02",X"10",X"02",X"12",X"05",X"12",X"06",X"15",X"05",X"15",X"06",X"17",X"06",
		X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"03",X"15",X"01",
		X"14",X"01",X"13",X"00",X"11",X"01",X"11",X"02",X"00",X"1D",X"00",X"1D",X"12",X"00",X"27",X"01",
		X"48",X"03",X"29",X"04",X"4A",X"03",X"4B",X"05",X"2C",X"04",X"2D",X"01",X"2D",X"07",X"2C",X"00",
		X"2C",X"02",X"2A",X"00",X"2A",X"02",X"48",X"08",X"29",X"06",X"28",X"01",X"29",X"01",X"29",X"00",
		X"29",X"06",X"29",X"01",X"2B",X"01",X"4C",X"03",X"2D",X"04",X"2F",X"03",X"30",X"09",X"2F",X"06",
		X"4D",X"07",X"2E",X"06",X"2C",X"02",X"49",X"07",X"4A",X"08",X"2B",X"06",X"28",X"00",X"28",X"02",
		X"27",X"00",X"28",X"01",X"29",X"01",X"2A",X"09",X"00",X"44",X"00",X"44",X"12",X"02",X"14",X"02",
		X"15",X"00",X"15",X"02",X"16",X"02",X"17",X"02",X"18",X"00",X"17",X"01",X"17",X"00",X"16",X"03",
		X"16",X"04",X"15",X"01",X"15",X"00",X"15",X"00",X"14",X"01",X"14",X"00",X"13",X"01",X"13",X"02",
		X"14",X"02",X"15",X"00",X"15",X"02",X"16",X"02",X"17",X"05",X"17",X"06",X"18",X"00",X"18",X"00",
		X"17",X"01",X"16",X"01",X"16",X"00",X"15",X"01",X"15",X"02",X"16",X"02",X"17",X"05",X"17",X"06",
		X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"17",X"00",X"16",X"01",X"14",X"01",X"12",X"03",
		X"12",X"04",X"12",X"02",X"13",X"02",X"14",X"05",X"14",X"06",X"17",X"02",X"18",X"00",X"17",X"01",
		X"17",X"00",X"17",X"00",X"16",X"03",X"16",X"04",X"15",X"01",X"14",X"01",X"14",X"00",X"14",X"02",
		X"15",X"05",X"15",X"06",X"17",X"05",X"17",X"06",X"18",X"00",X"17",X"03",X"17",X"04",X"16",X"01",
		X"15",X"01",X"13",X"01",X"00",X"44",X"00",X"44",X"29",X"02",X"28",X"02",X"27",X"02",X"47",X"03",
		X"28",X"04",X"29",X"01",X"4B",X"03",X"2C",X"04",X"2D",X"09",X"2C",X"06",X"2A",X"02",X"48",X"07",
		X"29",X"06",X"27",X"00",X"28",X"03",X"4A",X"03",X"2B",X"05",X"2C",X"09",X"2C",X"01",X"2D",X"09",
		X"2C",X"02",X"4A",X"07",X"2B",X"06",X"29",X"00",X"29",X"02",X"47",X"07",X"28",X"06",X"27",X"01",
		X"28",X"01",X"29",X"01",X"2A",X"01",X"2A",X"00",X"2A",X"02",X"29",X"00",X"29",X"02",X"28",X"02",
		X"27",X"07",X"27",X"04",X"48",X"03",X"29",X"05",X"4A",X"03",X"2B",X"04",X"2D",X"01",X"2E",X"09",
		X"2D",X"02",X"4B",X"07",X"2C",X"06",X"49",X"07",X"2A",X"06",X"28",X"02",X"28",X"01",X"29",X"01",
		X"2A",X"09",X"2A",X"01",X"2B",X"09",X"2A",X"02",X"29",X"02",X"28",X"02",X"28",X"04",X"49",X"03");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
