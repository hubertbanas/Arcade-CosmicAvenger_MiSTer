library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu3 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu3 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"60",X"FD",X"77",X"07",X"FD",X"36",X"08",X"00",X"DD",X"36",X"08",X"08",X"1E",X"09",X"CD",X"FB",
		X"06",X"C9",X"CD",X"7B",X"0B",X"FD",X"7E",X"14",X"E6",X"60",X"FE",X"40",X"CC",X"85",X"0B",X"DD",
		X"7E",X"02",X"FE",X"FD",X"38",X"23",X"C9",X"DD",X"7E",X"07",X"FE",X"0C",X"30",X"1B",X"A7",X"20",
		X"10",X"11",X"95",X"40",X"CD",X"21",X"07",X"1E",X"14",X"CD",X"0E",X"07",X"1E",X"02",X"CD",X"FB",
		X"06",X"CD",X"7B",X"0B",X"38",X"03",X"C3",X"C7",X"3D",X"DD",X"36",X"00",X"00",X"21",X"F8",X"63",
		X"35",X"C9",X"DD",X"34",X"09",X"DD",X"7E",X"05",X"FE",X"7C",X"38",X"0A",X"FE",X"8B",X"30",X"1B",
		X"DD",X"CB",X"09",X"76",X"20",X"15",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"11",X"80",X"00",X"19",
		X"DD",X"74",X"05",X"DD",X"75",X"06",X"DD",X"CB",X"09",X"B6",X"C9",X"DD",X"66",X"05",X"DD",X"6E",
		X"06",X"11",X"80",X"FF",X"19",X"DD",X"74",X"05",X"DD",X"75",X"06",X"DD",X"CB",X"09",X"F6",X"C9",
		X"00",X"01",X"00",X"00",X"01",X"00",X"DD",X"CB",X"00",X"66",X"C2",X"28",X"42",X"DD",X"7E",X"02",
		X"A7",X"28",X"0D",X"FA",X"C0",X"42",X"CD",X"7B",X"0B",X"D0",X"1E",X"0E",X"CD",X"FB",X"06",X"C9",
		X"DD",X"7E",X"05",X"C6",X"05",X"E6",X"F8",X"5F",X"CD",X"F6",X"0A",X"DD",X"86",X"03",X"C6",X"05",
		X"E6",X"F8",X"57",X"CD",X"03",X"0B",X"CD",X"15",X"0B",X"20",X"31",X"DD",X"7E",X"05",X"C6",X"09",
		X"E6",X"F8",X"5F",X"CD",X"F6",X"0A",X"DD",X"86",X"03",X"C6",X"09",X"E6",X"F8",X"57",X"CD",X"03",
		X"0B",X"CD",X"15",X"0B",X"20",X"2F",X"2A",X"7C",X"60",X"CB",X"3C",X"CB",X"1D",X"DD",X"56",X"05",
		X"DD",X"5E",X"06",X"19",X"DD",X"74",X"05",X"DD",X"75",X"06",X"18",X"46",X"ED",X"5B",X"7C",X"60",
		X"CB",X"3A",X"CB",X"1B",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"A7",X"ED",X"52",X"DD",X"74",X"05",
		X"DD",X"75",X"06",X"18",X"2D",X"DD",X"7E",X"05",X"4F",X"DD",X"96",X"0A",X"28",X"24",X"47",X"79",
		X"DD",X"96",X"0B",X"28",X"1D",X"30",X"02",X"ED",X"44",X"4F",X"78",X"CB",X"7F",X"28",X"02",X"ED",
		X"44",X"B9",X"30",X"08",X"DD",X"7E",X"0A",X"DD",X"77",X"05",X"18",X"06",X"DD",X"7E",X"0B",X"DD",
		X"77",X"05",X"ED",X"5B",X"7C",X"60",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"FD",X"7E",X"28",X"E6",
		X"1F",X"28",X"08",X"FE",X"04",X"30",X"04",X"CB",X"3A",X"CB",X"1B",X"CD",X"85",X"0B",X"30",X"06",
		X"1E",X"0E",X"CD",X"0E",X"07",X"C9",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"09",X"06",
		X"0E",X"0E",X"09",X"CD",X"41",X"0A",X"38",X"12",X"FD",X"21",X"60",X"63",X"CD",X"15",X"0A",X"28",
		X"12",X"06",X"17",X"0E",X"07",X"CD",X"41",X"0A",X"30",X"09",X"DD",X"CB",X"00",X"E6",X"FD",X"CB",
		X"00",X"E6",X"C9",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"5F",X"DD",X"7E",X"08",X"A7",
		X"28",X"13",X"DD",X"35",X"08",X"3A",X"E2",X"60",X"CB",X"2F",X"DD",X"BE",X"08",X"38",X"4C",X"DD",
		X"CB",X"00",X"86",X"18",X"46",X"CD",X"CB",X"42",X"20",X"41",X"3E",X"08",X"90",X"F6",X"80",X"77",
		X"E5",X"FD",X"E1",X"FD",X"36",X"02",X"00",X"DD",X"7E",X"03",X"D6",X"02",X"FD",X"77",X"03",X"DD",
		X"7E",X"04",X"FD",X"77",X"04",X"DD",X"7E",X"05",X"D6",X"03",X"FD",X"77",X"05",X"FD",X"36",X"06",
		X"00",X"FD",X"36",X"07",X"50",X"FD",X"36",X"08",X"00",X"CD",X"DA",X"42",X"DD",X"CB",X"00",X"C6",
		X"3A",X"E2",X"60",X"DD",X"77",X"08",X"1E",X"0B",X"CD",X"FB",X"06",X"06",X"C0",X"0E",X"50",X"16",
		X"04",X"3A",X"54",X"63",X"17",X"30",X"1D",X"DD",X"34",X"09",X"DD",X"CB",X"00",X"46",X"20",X"0A",
		X"DD",X"CB",X"09",X"5E",X"28",X"0E",X"0E",X"54",X"18",X"0A",X"0E",X"58",X"DD",X"CB",X"09",X"5E",
		X"28",X"02",X"0E",X"5C",X"CD",X"02",X"06",X"C9",X"DD",X"7E",X"07",X"FE",X"0C",X"D2",X"C0",X"42",
		X"A7",X"20",X"19",X"11",X"C7",X"42",X"DD",X"CB",X"00",X"46",X"20",X"03",X"11",X"CA",X"42",X"CD",
		X"21",X"07",X"1E",X"0E",X"CD",X"0E",X"07",X"1E",X"01",X"CD",X"FB",X"06",X"CD",X"7B",X"0B",X"38",
		X"6F",X"DD",X"7E",X"07",X"DD",X"34",X"07",X"E6",X"0C",X"28",X"06",X"FE",X"04",X"28",X"0B",X"18",
		X"42",X"01",X"98",X"C0",X"16",X"0D",X"CD",X"02",X"06",X"C9",X"11",X"F8",X"F8",X"CD",X"EF",X"0B",
		X"01",X"9C",X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",X"F8",X"08",X"CD",X"EF",X"0B",X"01",X"A0",
		X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",X"08",X"F8",X"CD",X"EF",X"0B",X"01",X"A4",X"C0",X"16",
		X"00",X"CD",X"08",X"06",X"11",X"08",X"08",X"CD",X"EF",X"0B",X"01",X"EC",X"C0",X"16",X"00",X"CD",
		X"08",X"06",X"C9",X"11",X"00",X"F8",X"CD",X"EF",X"0B",X"01",X"F0",X"C0",X"16",X"02",X"CD",X"08",
		X"06",X"11",X"00",X"08",X"CD",X"EF",X"0B",X"01",X"F4",X"C0",X"16",X"02",X"CD",X"08",X"06",X"C9",
		X"DD",X"36",X"00",X"00",X"C9",X"00",X"01",X"00",X"00",X"01",X"30",X"21",X"1C",X"65",X"11",X"0D",
		X"00",X"06",X"08",X"CB",X"7E",X"C8",X"19",X"10",X"FA",X"C9",X"3A",X"57",X"63",X"DD",X"96",X"03",
		X"30",X"02",X"ED",X"44",X"47",X"3A",X"59",X"63",X"DD",X"96",X"05",X"30",X"02",X"ED",X"44",X"4F",
		X"B8",X"30",X"1D",X"69",X"59",X"26",X"00",X"16",X"00",X"29",X"29",X"19",X"58",X"ED",X"52",X"38",
		X"2C",X"69",X"59",X"26",X"00",X"29",X"19",X"EB",X"68",X"29",X"ED",X"52",X"38",X"31",X"18",X"26",
		X"68",X"58",X"26",X"00",X"16",X"00",X"29",X"29",X"19",X"59",X"ED",X"52",X"38",X"33",X"68",X"58",
		X"26",X"00",X"29",X"19",X"EB",X"69",X"29",X"ED",X"52",X"38",X"14",X"18",X"1B",X"ED",X"5B",X"80",
		X"43",X"2A",X"82",X"43",X"18",X"22",X"ED",X"5B",X"84",X"43",X"2A",X"86",X"43",X"18",X"19",X"ED",
		X"5B",X"88",X"43",X"2A",X"8A",X"43",X"18",X"10",X"ED",X"5B",X"8C",X"43",X"2A",X"8E",X"43",X"18",
		X"07",X"ED",X"5B",X"90",X"43",X"2A",X"92",X"43",X"3A",X"59",X"63",X"DD",X"96",X"05",X"DC",X"78",
		X"43",X"FD",X"74",X"0B",X"FD",X"75",X"0C",X"EB",X"3A",X"57",X"63",X"DD",X"96",X"03",X"DC",X"78",
		X"43",X"FD",X"74",X"09",X"FD",X"75",X"0A",X"C9",X"7D",X"2F",X"6F",X"7C",X"2F",X"67",X"23",X"C9",
		X"00",X"03",X"00",X"00",X"C6",X"02",X"26",X"01",X"1F",X"02",X"1F",X"02",X"26",X"01",X"C6",X"02",
		X"00",X"00",X"00",X"03",X"DD",X"CB",X"00",X"5E",X"C2",X"8B",X"45",X"DD",X"CB",X"00",X"66",X"C2",
		X"68",X"44",X"CD",X"7B",X"0B",X"DA",X"82",X"45",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"DD",X"CB",
		X"00",X"6E",X"20",X"0F",X"11",X"80",X"00",X"19",X"7C",X"FE",X"8A",X"38",X"15",X"DD",X"CB",X"00",
		X"EE",X"18",X"15",X"11",X"80",X"FF",X"19",X"7C",X"FE",X"7C",X"30",X"06",X"DD",X"CB",X"00",X"AE",
		X"18",X"06",X"DD",X"74",X"05",X"DD",X"75",X"06",X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",
		X"C2",X"5E",X"44",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"09",X"06",X"0C",X"0E",X"08",
		X"CD",X"41",X"0A",X"38",X"60",X"FD",X"21",X"60",X"63",X"CD",X"15",X"0A",X"28",X"09",X"06",X"15",
		X"0E",X"06",X"CD",X"41",X"0A",X"38",X"4E",X"FD",X"21",X"68",X"63",X"CD",X"15",X"0A",X"28",X"0F",
		X"FD",X"CB",X"00",X"46",X"20",X"09",X"06",X"08",X"0E",X"06",X"CD",X"41",X"0A",X"38",X"36",X"FD",
		X"21",X"79",X"63",X"CD",X"15",X"0A",X"28",X"0F",X"FD",X"CB",X"00",X"46",X"20",X"09",X"06",X"08",
		X"0E",X"06",X"CD",X"41",X"0A",X"38",X"1E",X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"06",X"0D",
		X"0E",X"09",X"26",X"08",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"07",X"FD",X"19",
		X"25",X"20",X"F1",X"18",X"09",X"DD",X"CB",X"00",X"E6",X"FD",X"CB",X"00",X"E6",X"C9",X"06",X"C0",
		X"0E",X"60",X"16",X"0C",X"CD",X"02",X"06",X"C9",X"DD",X"7E",X"07",X"FE",X"28",X"D2",X"82",X"45",
		X"A7",X"20",X"0B",X"11",X"48",X"46",X"CD",X"21",X"07",X"1E",X"11",X"CD",X"FB",X"06",X"CD",X"7B",
		X"0B",X"DA",X"82",X"45",X"DD",X"7E",X"07",X"CD",X"A9",X"0B",X"3A",X"03",X"60",X"DD",X"AE",X"00",
		X"E6",X"03",X"C2",X"7E",X"45",X"DD",X"7E",X"07",X"CD",X"1F",X"0A",X"FD",X"21",X"54",X"63",X"CD",
		X"15",X"0A",X"28",X"0A",X"06",X"07",X"0E",X"03",X"CD",X"39",X"0A",X"DA",X"7A",X"45",X"FD",X"21",
		X"60",X"63",X"CD",X"15",X"0A",X"28",X"0A",X"06",X"10",X"0E",X"01",X"CD",X"39",X"0A",X"DA",X"7A",
		X"45",X"FD",X"21",X"68",X"63",X"CD",X"15",X"0A",X"28",X"10",X"FD",X"CB",X"00",X"46",X"20",X"0A",
		X"06",X"03",X"0E",X"01",X"CD",X"39",X"0A",X"DA",X"7A",X"45",X"FD",X"21",X"79",X"63",X"CD",X"15",
		X"0A",X"28",X"10",X"FD",X"CB",X"00",X"46",X"20",X"0A",X"06",X"03",X"0E",X"01",X"CD",X"39",X"0A",
		X"DA",X"7A",X"45",X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",X"06",X"0C",X"CD",X"15",X"0A",X"28",
		X"0B",X"C5",X"06",X"08",X"0E",X"08",X"CD",X"39",X"0A",X"C1",X"38",X"6E",X"FD",X"19",X"10",X"EC",
		X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"06",X"08",X"CD",X"15",X"0A",X"28",X"0B",X"C5",X"06",
		X"08",X"0E",X"04",X"CD",X"39",X"0A",X"C1",X"38",X"51",X"FD",X"19",X"10",X"EC",X"FD",X"21",X"DC",
		X"64",X"11",X"08",X"00",X"06",X"08",X"CD",X"15",X"0A",X"28",X"15",X"C5",X"06",X"05",X"0E",X"05",
		X"FD",X"CB",X"00",X"5E",X"28",X"04",X"06",X"04",X"0E",X"06",X"CD",X"39",X"0A",X"C1",X"38",X"2A",
		X"FD",X"19",X"10",X"E2",X"FD",X"21",X"1C",X"65",X"11",X"0D",X"00",X"06",X"08",X"CD",X"15",X"0A",
		X"28",X"12",X"C5",X"D5",X"01",X"00",X"00",X"FD",X"7E",X"07",X"CD",X"0E",X"4C",X"CD",X"39",X"0A",
		X"D1",X"C1",X"38",X"06",X"FD",X"19",X"10",X"E5",X"18",X"04",X"FD",X"CB",X"00",X"E6",X"DD",X"34",
		X"07",X"C9",X"DD",X"36",X"00",X"00",X"21",X"F6",X"63",X"35",X"C9",X"DD",X"CB",X"00",X"66",X"C2",
		X"35",X"46",X"CD",X"7B",X"0B",X"38",X"EB",X"21",X"00",X"01",X"DD",X"56",X"05",X"DD",X"5E",X"06",
		X"19",X"DD",X"74",X"05",X"DD",X"75",X"06",X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"C2",
		X"2B",X"46",X"06",X"04",X"0E",X"06",X"CD",X"60",X"0A",X"28",X"09",X"DD",X"CB",X"00",X"EE",X"DD",
		X"CB",X"00",X"E6",X"C9",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"09",X"06",X"0B",X"0E",
		X"09",X"CD",X"41",X"0A",X"38",X"4C",X"FD",X"21",X"60",X"63",X"CD",X"15",X"0A",X"28",X"09",X"06",
		X"14",X"0E",X"07",X"CD",X"41",X"0A",X"38",X"3A",X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",X"26",
		X"0C",X"06",X"0C",X"0E",X"0E",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"23",X"FD",
		X"19",X"25",X"20",X"F1",X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"26",X"08",X"06",X"0C",X"0E",
		X"0A",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"07",X"FD",X"19",X"25",X"20",X"F1",
		X"18",X"09",X"DD",X"CB",X"00",X"E6",X"FD",X"CB",X"00",X"E6",X"C9",X"06",X"C0",X"0E",X"64",X"16",
		X"03",X"CD",X"02",X"06",X"C9",X"DD",X"CB",X"00",X"6E",X"CA",X"68",X"44",X"DD",X"7E",X"07",X"A7",
		X"C2",X"68",X"44",X"C3",X"79",X"44",X"00",X"00",X"50",X"00",X"00",X"50",X"DD",X"CB",X"00",X"66",
		X"C2",X"9F",X"4A",X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"C2",X"03",X"47",X"FD",X"21",
		X"54",X"63",X"CD",X"15",X"0A",X"28",X"0F",X"01",X"03",X"07",X"DD",X"7E",X"07",X"CD",X"0E",X"4C",
		X"CD",X"41",X"0A",X"DA",X"FA",X"46",X"FD",X"21",X"60",X"63",X"CD",X"15",X"0A",X"28",X"0E",X"01",
		X"01",X"10",X"DD",X"7E",X"07",X"CD",X"0E",X"4C",X"CD",X"41",X"0A",X"38",X"6D",X"FD",X"21",X"68",
		X"63",X"CD",X"15",X"0A",X"28",X"0E",X"01",X"02",X"03",X"DD",X"7E",X"07",X"CD",X"0E",X"4C",X"CD",
		X"41",X"0A",X"38",X"56",X"FD",X"21",X"79",X"63",X"CD",X"15",X"0A",X"28",X"0E",X"01",X"02",X"03",
		X"DD",X"7E",X"07",X"CD",X"0E",X"4C",X"CD",X"41",X"0A",X"38",X"3F",X"DD",X"7E",X"00",X"E6",X"07",
		X"28",X"41",X"FD",X"21",X"6A",X"65",X"11",X"F3",X"FF",X"47",X"D6",X"07",X"28",X"07",X"ED",X"44",
		X"FD",X"19",X"3D",X"20",X"FB",X"D9",X"01",X"00",X"00",X"DD",X"7E",X"07",X"CD",X"0E",X"4C",X"D9",
		X"CD",X"15",X"0A",X"28",X"0F",X"D9",X"C5",X"FD",X"7E",X"07",X"CD",X"0E",X"4C",X"CD",X"41",X"0A",
		X"C1",X"D9",X"38",X"06",X"FD",X"19",X"10",X"E8",X"18",X"09",X"DD",X"CB",X"00",X"E6",X"FD",X"CB",
		X"00",X"E6",X"C9",X"DD",X"7E",X"07",X"E6",X"70",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"17",
		X"47",X"19",X"5E",X"23",X"56",X"EB",X"E9",X"27",X"47",X"80",X"47",X"EC",X"47",X"CC",X"48",X"88",
		X"49",X"EA",X"49",X"39",X"4A",X"C8",X"4B",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"ED",X"5B",X"E3",
		X"60",X"A7",X"ED",X"52",X"7C",X"FE",X"40",X"38",X"44",X"DD",X"74",X"05",X"DD",X"75",X"06",X"CD",
		X"7B",X"0B",X"38",X"39",X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"20",X"1C",X"FD",X"21",
		X"80",X"64",X"11",X"0A",X"00",X"26",X"08",X"06",X"0C",X"0E",X"0A",X"CD",X"15",X"0A",X"28",X"05",
		X"CD",X"41",X"0A",X"38",X"0F",X"FD",X"19",X"25",X"20",X"F1",X"06",X"C0",X"0E",X"14",X"16",X"06",
		X"CD",X"02",X"06",X"C9",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"E6",X"C9",X"C3",X"C8",X"4B",
		X"CD",X"7B",X"0B",X"38",X"64",X"DD",X"CB",X"09",X"66",X"20",X"05",X"DD",X"34",X"09",X"18",X"08",
		X"3A",X"59",X"63",X"DD",X"BE",X"05",X"30",X"4C",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"ED",X"5B",
		X"E3",X"60",X"A7",X"ED",X"52",X"7C",X"FE",X"44",X"38",X"3A",X"DD",X"74",X"05",X"DD",X"75",X"06",
		X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"20",X"1C",X"FD",X"21",X"80",X"64",X"11",X"0A",
		X"00",X"26",X"08",X"06",X"0A",X"0E",X"08",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",
		X"0F",X"FD",X"19",X"25",X"20",X"F1",X"06",X"80",X"0E",X"6F",X"16",X"0C",X"CD",X"02",X"06",X"C9",
		X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"E6",X"C9",X"C3",X"C8",X"4B",X"DD",X"CB",X"00",X"5E",
		X"20",X"0F",X"CD",X"B6",X"48",X"3A",X"59",X"63",X"BC",X"38",X"7B",X"DD",X"CB",X"00",X"DE",X"18",
		X"75",X"ED",X"5B",X"7C",X"60",X"21",X"C0",X"03",X"A7",X"ED",X"52",X"DD",X"56",X"03",X"DD",X"5E",
		X"04",X"19",X"7C",X"FE",X"F8",X"D2",X"C8",X"4B",X"FE",X"08",X"38",X"06",X"DD",X"74",X"03",X"DD",
		X"75",X"04",X"DD",X"34",X"09",X"DD",X"7E",X"09",X"E6",X"01",X"20",X"12",X"3A",X"59",X"63",X"DD",
		X"BE",X"05",X"28",X"0A",X"30",X"05",X"CD",X"B6",X"48",X"18",X"03",X"CD",X"BB",X"48",X"3A",X"03",
		X"60",X"DD",X"AE",X"00",X"E6",X"03",X"20",X"53",X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",X"26",
		X"0C",X"06",X"0F",X"0E",X"0C",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"4E",X"FD",
		X"19",X"25",X"20",X"F1",X"FD",X"21",X"D0",X"64",X"CD",X"15",X"0A",X"28",X"09",X"06",X"0E",X"0E",
		X"0A",X"CD",X"41",X"0A",X"38",X"37",X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"26",X"08",X"06",
		X"0F",X"0E",X"08",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"20",X"FD",X"19",X"25",
		X"20",X"F1",X"06",X"07",X"0E",X"04",X"CD",X"60",X"0A",X"20",X"16",X"06",X"C0",X"0E",X"28",X"16",
		X"03",X"DD",X"CB",X"00",X"5E",X"28",X"02",X"0E",X"2C",X"CD",X"02",X"06",X"C9",X"FD",X"CB",X"00",
		X"E6",X"DD",X"CB",X"00",X"E6",X"C9",X"11",X"00",X"FF",X"18",X"03",X"11",X"00",X"01",X"DD",X"66",
		X"05",X"DD",X"6E",X"06",X"19",X"DD",X"74",X"05",X"DD",X"75",X"06",X"C9",X"DD",X"CB",X"00",X"5E",
		X"20",X"30",X"2A",X"7C",X"60",X"11",X"00",X"02",X"19",X"EB",X"DD",X"66",X"03",X"DD",X"6E",X"04",
		X"CD",X"85",X"0B",X"DA",X"85",X"49",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"11",X"00",X"02",X"19",
		X"DD",X"74",X"05",X"DD",X"75",X"06",X"7C",X"DD",X"BE",X"09",X"38",X"1A",X"DD",X"CB",X"00",X"DE",
		X"18",X"14",X"2A",X"7C",X"60",X"ED",X"5B",X"E5",X"60",X"19",X"EB",X"DD",X"66",X"03",X"DD",X"6E",
		X"04",X"CD",X"85",X"0B",X"38",X"6F",X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"20",X"4A",
		X"01",X"03",X"08",X"CD",X"60",X"0A",X"20",X"58",X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"26",
		X"08",X"06",X"10",X"0E",X"07",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"3D",X"FD",
		X"19",X"25",X"20",X"F1",X"FD",X"21",X"DC",X"64",X"11",X"08",X"00",X"26",X"08",X"CD",X"15",X"0A",
		X"28",X"13",X"06",X"0D",X"0E",X"08",X"FD",X"CB",X"00",X"5E",X"28",X"04",X"06",X"0C",X"0E",X"09",
		X"CD",X"41",X"0A",X"38",X"17",X"FD",X"19",X"25",X"20",X"E3",X"06",X"F0",X"0E",X"28",X"16",X"03",
		X"DD",X"CB",X"00",X"5E",X"28",X"02",X"0E",X"2C",X"CD",X"02",X"06",X"C9",X"FD",X"CB",X"00",X"E6",
		X"DD",X"CB",X"00",X"E6",X"C9",X"C3",X"C8",X"4B",X"CD",X"D2",X"4B",X"DA",X"C8",X"4B",X"3A",X"03",
		X"60",X"DD",X"AE",X"00",X"E6",X"03",X"20",X"37",X"06",X"01",X"0E",X"00",X"CD",X"60",X"0A",X"20",
		X"44",X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",X"26",X"0C",X"06",X"09",X"0E",X"08",X"CD",X"15",
		X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"29",X"FD",X"19",X"25",X"20",X"F1",X"FD",X"21",X"D0",
		X"64",X"CD",X"15",X"0A",X"28",X"09",X"06",X"08",X"0E",X"06",X"CD",X"41",X"0A",X"38",X"12",X"06",
		X"80",X"DD",X"CB",X"09",X"7E",X"28",X"02",X"CB",X"E8",X"0E",X"72",X"16",X"0D",X"CD",X"02",X"06",
		X"C9",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"E6",X"C9",X"CD",X"D2",X"4B",X"38",X"42",X"3A",
		X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"20",X"25",X"06",X"04",X"0E",X"03",X"CD",X"60",X"0A",
		X"20",X"2A",X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"26",X"08",X"06",X"0C",X"0E",X"07",X"CD",
		X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"0F",X"FD",X"19",X"25",X"20",X"F1",X"06",X"80",
		X"0E",X"71",X"16",X"02",X"CD",X"02",X"06",X"C9",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"E6",
		X"C9",X"1E",X"0B",X"CD",X"0E",X"07",X"C3",X"C8",X"4B",X"2A",X"7C",X"60",X"11",X"00",X"03",X"19",
		X"EB",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"CD",X"85",X"0B",X"38",X"4B",X"3A",X"03",X"60",X"DD",
		X"AE",X"00",X"E6",X"03",X"20",X"2E",X"01",X"02",X"04",X"CD",X"60",X"0A",X"20",X"34",X"FD",X"21",
		X"DC",X"64",X"11",X"08",X"00",X"26",X"08",X"CD",X"15",X"0A",X"28",X"13",X"06",X"09",X"0E",X"07",
		X"FD",X"CB",X"00",X"5E",X"28",X"04",X"06",X"08",X"0E",X"08",X"CD",X"41",X"0A",X"38",X"0F",X"FD",
		X"19",X"25",X"20",X"E3",X"06",X"80",X"0E",X"73",X"16",X"0C",X"CD",X"02",X"06",X"C9",X"FD",X"CB",
		X"00",X"E6",X"DD",X"CB",X"00",X"E6",X"C9",X"1E",X"09",X"CD",X"0E",X"07",X"C3",X"C8",X"4B",X"DD",
		X"7E",X"07",X"E6",X"70",X"FE",X"10",X"28",X"51",X"DD",X"7E",X"08",X"FE",X"0C",X"30",X"47",X"A7",
		X"20",X"32",X"DD",X"7E",X"07",X"E6",X"70",X"0F",X"0F",X"0F",X"47",X"0F",X"80",X"5F",X"16",X"00",
		X"21",X"34",X"4C",X"19",X"EB",X"CD",X"21",X"07",X"DD",X"7E",X"07",X"E6",X"07",X"FE",X"05",X"38",
		X"0E",X"20",X"07",X"1E",X"0B",X"CD",X"0E",X"07",X"18",X"05",X"1E",X"09",X"CD",X"0E",X"07",X"1E",
		X"12",X"CD",X"FB",X"06",X"CD",X"7B",X"0B",X"38",X"0D",X"DD",X"7E",X"08",X"21",X"A3",X"0B",X"CD",
		X"93",X"0B",X"DD",X"34",X"08",X"C9",X"C3",X"C8",X"4B",X"DD",X"7E",X"08",X"FE",X"28",X"D2",X"C8",
		X"4B",X"A7",X"20",X"05",X"1E",X"11",X"CD",X"FB",X"06",X"CD",X"7B",X"0B",X"DA",X"C8",X"4B",X"DD",
		X"7E",X"08",X"CD",X"A9",X"0B",X"3A",X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"C2",X"C4",X"4B",
		X"DD",X"7E",X"08",X"CD",X"1F",X"0A",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"0A",X"06",
		X"07",X"0E",X"03",X"CD",X"39",X"0A",X"DA",X"C0",X"4B",X"FD",X"21",X"60",X"63",X"CD",X"15",X"0A",
		X"28",X"09",X"06",X"10",X"0E",X"01",X"CD",X"39",X"0A",X"38",X"75",X"FD",X"21",X"68",X"63",X"CD",
		X"15",X"0A",X"28",X"0F",X"FD",X"CB",X"00",X"46",X"20",X"09",X"06",X"03",X"0E",X"01",X"CD",X"39",
		X"0A",X"38",X"5D",X"FD",X"21",X"79",X"63",X"CD",X"15",X"0A",X"28",X"0F",X"FD",X"CB",X"00",X"46",
		X"20",X"09",X"06",X"03",X"0E",X"01",X"CD",X"39",X"0A",X"38",X"45",X"FD",X"21",X"80",X"64",X"11",
		X"0A",X"00",X"06",X"08",X"CD",X"15",X"0A",X"28",X"0B",X"C5",X"06",X"08",X"0E",X"04",X"CD",X"39",
		X"0A",X"C1",X"38",X"2C",X"FD",X"19",X"10",X"EC",X"FD",X"21",X"1C",X"65",X"D9",X"11",X"0D",X"00",
		X"06",X"08",X"CD",X"15",X"0A",X"28",X"12",X"D9",X"01",X"00",X"00",X"FD",X"7E",X"07",X"E5",X"CD",
		X"0E",X"4C",X"E1",X"CD",X"39",X"0A",X"38",X"08",X"D9",X"FD",X"19",X"10",X"E5",X"D9",X"18",X"04",
		X"FD",X"CB",X"00",X"E6",X"DD",X"34",X"08",X"C9",X"DD",X"36",X"00",X"00",X"21",X"01",X"60",X"CB",
		X"FE",X"C9",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"DD",X"66",X"09",X"DD",X"6E",X"0A",X"19",X"7C",
		X"FE",X"08",X"38",X"28",X"FE",X"F8",X"30",X"24",X"DD",X"74",X"03",X"DD",X"75",X"04",X"DD",X"56",
		X"05",X"DD",X"5E",X"06",X"DD",X"66",X"0B",X"DD",X"6E",X"0C",X"19",X"7C",X"FE",X"40",X"38",X"0C",
		X"FE",X"C0",X"30",X"08",X"DD",X"74",X"05",X"DD",X"75",X"06",X"A7",X"C9",X"37",X"C9",X"E6",X"70",
		X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"22",X"4C",X"19",X"7E",X"80",X"47",X"23",X"7E",X"81",
		X"4F",X"C9",X"04",X"08",X"02",X"04",X"07",X"04",X"08",X"03",X"01",X"00",X"04",X"03",X"04",X"02",
		X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"00",X"00",X"00",X"30",X"00",X"00",X"30",X"00",X"00",
		X"50",X"00",X"00",X"30",X"00",X"00",X"50",X"00",X"00",X"00",X"EF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"34",X"50",X"39",X"50",X"3E",X"50",X"43",X"50",X"48",X"50",X"4B",X"50",X"4E",X"50",X"50",X"50",
		X"52",X"50",X"54",X"50",X"57",X"50",X"5A",X"50",X"62",X"50",X"5F",X"50",X"5C",X"50",X"65",X"50",
		X"67",X"50",X"6A",X"50",X"6D",X"50",X"70",X"50",X"73",X"50",X"76",X"50",X"79",X"50",X"7C",X"50",
		X"82",X"50",X"88",X"50",X"04",X"20",X"30",X"60",X"70",X"04",X"20",X"30",X"60",X"70",X"04",X"20",
		X"30",X"60",X"70",X"04",X"20",X"30",X"60",X"70",X"02",X"60",X"70",X"02",X"40",X"50",X"01",X"00",
		X"01",X"00",X"01",X"00",X"02",X"20",X"30",X"02",X"00",X"10",X"01",X"00",X"02",X"20",X"30",X"02",
		X"20",X"30",X"02",X"00",X"10",X"01",X"00",X"02",X"00",X"10",X"02",X"00",X"10",X"02",X"20",X"30",
		X"02",X"00",X"10",X"02",X"00",X"10",X"02",X"00",X"10",X"02",X"00",X"10",X"FF",X"9A",X"5C",X"03",
		X"0C",X"5D",X"FF",X"51",X"5D",X"03",X"9D",X"5D",X"02",X"20",X"30",X"FD",X"21",X"00",X"6C",X"DD",
		X"21",X"06",X"6C",X"FD",X"36",X"02",X"00",X"01",X"00",X"1A",X"21",X"29",X"52",X"DD",X"7E",X"00",
		X"E6",X"03",X"20",X"07",X"DD",X"36",X"00",X"00",X"C3",X"04",X"52",X"E5",X"DD",X"CB",X"00",X"56",
		X"28",X"15",X"DD",X"36",X"00",X"00",X"CF",X"23",X"36",X"00",X"FD",X"7E",X"02",X"A7",X"C2",X"03",
		X"52",X"CD",X"91",X"52",X"C3",X"03",X"52",X"FD",X"34",X"02",X"CB",X"47",X"28",X"1B",X"DD",X"CB",
		X"00",X"86",X"DD",X"CB",X"00",X"CE",X"CF",X"71",X"23",X"36",X"80",X"FD",X"7E",X"02",X"FE",X"01",
		X"C2",X"03",X"52",X"CD",X"91",X"52",X"C3",X"03",X"52",X"C5",X"DD",X"E5",X"CF",X"E5",X"DD",X"E1",
		X"DD",X"CB",X"01",X"76",X"28",X"09",X"DD",X"35",X"02",X"20",X"0F",X"DD",X"CB",X"01",X"B6",X"EB",
		X"CF",X"FD",X"E5",X"01",X"08",X"51",X"C5",X"E9",X"FD",X"E1",X"FD",X"7E",X"02",X"FE",X"01",X"C2",
		X"00",X"52",X"DD",X"CB",X"01",X"7E",X"CA",X"00",X"52",X"DD",X"6E",X"00",X"26",X"00",X"29",X"11",
		X"00",X"50",X"19",X"CF",X"7E",X"FE",X"FF",X"CA",X"87",X"51",X"47",X"23",X"7E",X"23",X"E5",X"21",
		X"00",X"B0",X"FE",X"40",X"38",X"05",X"D6",X"40",X"21",X"00",X"C0",X"87",X"C6",X"80",X"4F",X"FE",
		X"E0",X"28",X"1E",X"DD",X"7E",X"03",X"E6",X"0F",X"81",X"77",X"DD",X"7E",X"03",X"E6",X"F0",X"0F",
		X"0F",X"0F",X"0F",X"5F",X"DD",X"7E",X"04",X"E6",X"03",X"07",X"07",X"07",X"07",X"83",X"77",X"18",
		X"11",X"DD",X"CB",X"04",X"7E",X"28",X"0B",X"DD",X"CB",X"04",X"BE",X"DD",X"7E",X"03",X"E6",X"07",
		X"81",X"77",X"DD",X"7E",X"05",X"2F",X"E6",X"0F",X"81",X"C6",X"10",X"77",X"E1",X"11",X"03",X"00",
		X"DD",X"19",X"10",X"A8",X"C3",X"00",X"52",X"FD",X"36",X"03",X"02",X"21",X"00",X"B0",X"FD",X"36",
		X"04",X"03",X"01",X"80",X"90",X"DD",X"7E",X"04",X"2F",X"E6",X"0F",X"80",X"47",X"DD",X"23",X"DD",
		X"7E",X"04",X"A7",X"20",X"06",X"78",X"F6",X"0F",X"77",X"18",X"23",X"E5",X"6F",X"26",X"00",X"29",
		X"11",X"D5",X"52",X"19",X"CF",X"7D",X"E6",X"0F",X"81",X"57",X"7D",X"E6",X"F0",X"0F",X"0F",X"0F",
		X"0F",X"6F",X"7C",X"E6",X"03",X"07",X"07",X"07",X"07",X"85",X"E1",X"72",X"77",X"70",X"E5",X"21",
		X"20",X"20",X"09",X"44",X"4D",X"E1",X"DD",X"23",X"FD",X"35",X"04",X"20",X"C2",X"DD",X"7E",X"04",
		X"DD",X"CB",X"04",X"BE",X"CB",X"77",X"20",X"04",X"06",X"FF",X"18",X"08",X"CB",X"7F",X"28",X"04",
		X"E6",X"07",X"81",X"77",X"70",X"DD",X"23",X"FD",X"35",X"03",X"21",X"00",X"C0",X"C2",X"8E",X"51",
		X"DD",X"E1",X"C1",X"E1",X"11",X"04",X"00",X"19",X"DD",X"23",X"0C",X"79",X"FE",X"06",X"20",X"0A",
		X"FD",X"7E",X"02",X"FD",X"77",X"05",X"FD",X"36",X"02",X"00",X"05",X"C2",X"9D",X"50",X"FD",X"7E",
		X"02",X"FD",X"86",X"05",X"C0",X"CD",X"91",X"52",X"C9",X"20",X"6C",X"26",X"58",X"39",X"6C",X"26",
		X"58",X"52",X"6C",X"26",X"58",X"6B",X"6C",X"26",X"58",X"84",X"6C",X"A4",X"58",X"8F",X"6C",X"C4",
		X"58",X"99",X"6C",X"07",X"59",X"A1",X"6C",X"07",X"59",X"A9",X"6C",X"22",X"59",X"B6",X"6C",X"76",
		X"59",X"C0",X"6C",X"AB",X"59",X"CE",X"6C",X"22",X"59",X"F1",X"6C",X"15",X"5A",X"E6",X"6C",X"A4",
		X"58",X"DB",X"6C",X"A4",X"58",X"02",X"6D",X"07",X"59",X"0A",X"6D",X"7F",X"5A",X"1B",X"6D",X"06",
		X"5B",X"26",X"6D",X"79",X"5B",X"30",X"6D",X"7F",X"5A",X"41",X"6D",X"AD",X"5B",X"51",X"6D",X"7F",
		X"5A",X"62",X"6D",X"62",X"5C",X"6E",X"6D",X"3D",X"53",X"CE",X"6D",X"3D",X"53",X"2E",X"6E",X"A4",
		X"58",X"3E",X"9F",X"32",X"00",X"B0",X"32",X"00",X"C0",X"C6",X"20",X"30",X"F6",X"C9",X"DD",X"36",
		X"01",X"00",X"DD",X"5E",X"00",X"16",X"00",X"21",X"06",X"6C",X"19",X"36",X"00",X"3A",X"02",X"6C",
		X"FE",X"01",X"C0",X"CD",X"91",X"52",X"C9",X"00",X"01",X"80",X"01",X"00",X"02",X"00",X"03",X"00",
		X"04",X"00",X"06",X"00",X"08",X"00",X"0C",X"00",X"10",X"00",X"18",X"00",X"20",X"AA",X"00",X"55",
		X"01",X"AA",X"02",X"55",X"05",X"00",X"00",X"F8",X"03",X"BF",X"03",X"89",X"03",X"56",X"03",X"26",
		X"03",X"FA",X"02",X"CE",X"02",X"A6",X"02",X"80",X"02",X"5C",X"02",X"3A",X"02",X"1A",X"02",X"FC",
		X"01",X"DF",X"01",X"C4",X"01",X"AB",X"01",X"93",X"01",X"7D",X"01",X"67",X"01",X"53",X"01",X"40",
		X"01",X"2E",X"01",X"1D",X"01",X"0D",X"01",X"FE",X"00",X"F0",X"00",X"E2",X"00",X"D6",X"00",X"CA",
		X"00",X"BE",X"00",X"B4",X"00",X"AA",X"00",X"A0",X"00",X"97",X"00",X"8F",X"00",X"87",X"00",X"7F",
		X"00",X"78",X"00",X"71",X"00",X"6B",X"00",X"65",X"00",X"5F",X"00",X"5A",X"00",X"55",X"00",X"50",
		X"00",X"4B",X"00",X"47",X"00",X"43",X"00",X"3F",X"00",X"3C",X"00",X"39",X"00",X"DD",X"CB",X"01",
		X"6E",X"20",X"5B",X"DD",X"E5",X"E1",X"23",X"23",X"AF",X"01",X"01",X"5E",X"D7",X"DD",X"CB",X"01",
		X"EE",X"DD",X"5E",X"00",X"CB",X"23",X"16",X"00",X"21",X"00",X"50",X"19",X"CF",X"23",X"CF",X"DD",
		X"E5",X"FD",X"E1",X"01",X"0E",X"00",X"FD",X"09",X"FD",X"CB",X"00",X"FE",X"46",X"23",X"4E",X"23",
		X"FD",X"75",X"0A",X"FD",X"74",X"0B",X"FD",X"71",X"0C",X"FD",X"70",X"0D",X"1A",X"DD",X"77",X"03",
		X"FE",X"01",X"C8",X"13",X"EB",X"CF",X"11",X"29",X"00",X"FD",X"19",X"FD",X"CB",X"00",X"FE",X"4E",
		X"23",X"FD",X"75",X"0A",X"FD",X"74",X"0B",X"FD",X"71",X"0C",X"FD",X"70",X"0D",X"C9",X"DD",X"7E",
		X"03",X"A7",X"20",X"04",X"CD",X"9E",X"52",X"C9",X"DD",X"CB",X"03",X"46",X"28",X"23",X"DD",X"E5",
		X"11",X"0E",X"00",X"DD",X"19",X"DD",X"E5",X"FD",X"E1",X"DD",X"E1",X"DD",X"E5",X"11",X"04",X"00",
		X"DD",X"19",X"CD",X"F9",X"53",X"DD",X"E1",X"FD",X"CB",X"00",X"7E",X"20",X"04",X"DD",X"CB",X"03",
		X"86",X"DD",X"CB",X"03",X"4E",X"C8",X"DD",X"E5",X"11",X"37",X"00",X"DD",X"19",X"DD",X"E5",X"FD",
		X"E1",X"DD",X"E1",X"DD",X"E5",X"11",X"09",X"00",X"DD",X"19",X"CD",X"F9",X"53",X"DD",X"E1",X"FD",
		X"CB",X"00",X"7E",X"C0",X"DD",X"CB",X"03",X"8E",X"C9",X"06",X"05",X"21",X"2C",X"54",X"FD",X"E5",
		X"FD",X"CB",X"00",X"7E",X"28",X"1B",X"FD",X"CB",X"00",X"76",X"28",X"09",X"FD",X"35",X"01",X"20",
		X"10",X"FD",X"CB",X"00",X"B6",X"C5",X"CF",X"D5",X"11",X"1D",X"54",X"D5",X"E9",X"E1",X"C1",X"18",
		X"02",X"23",X"23",X"FD",X"23",X"FD",X"23",X"10",X"D7",X"FD",X"E1",X"C9",X"36",X"54",X"3B",X"56",
		X"79",X"56",X"82",X"56",X"AB",X"56",X"CD",X"B0",X"55",X"CB",X"7C",X"20",X"07",X"CB",X"6D",X"C2",
		X"21",X"55",X"18",X"38",X"FD",X"36",X"06",X"00",X"DD",X"36",X"00",X"00",X"DD",X"36",X"01",X"00",
		X"DD",X"36",X"02",X"00",X"DD",X"36",X"03",X"00",X"DD",X"36",X"04",X"00",X"7C",X"E6",X"70",X"0F",
		X"0F",X"0F",X"5F",X"16",X"00",X"21",X"6C",X"54",X"19",X"CF",X"E9",X"C9",X"6B",X"54",X"35",X"55",
		X"4A",X"55",X"60",X"55",X"6B",X"54",X"6B",X"54",X"6B",X"54",X"AB",X"55",X"FD",X"7E",X"10",X"A7",
		X"20",X"18",X"FD",X"36",X"06",X"00",X"DD",X"36",X"01",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",
		X"03",X"00",X"FD",X"7E",X"0C",X"E6",X"0F",X"DD",X"77",X"00",X"CB",X"74",X"C2",X"00",X"55",X"7D",
		X"E6",X"0F",X"CD",X"D9",X"55",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"F6",X"FD",X"7E",X"0F",X"E6",
		X"3F",X"20",X"05",X"DD",X"36",X"00",X"00",X"C9",X"FD",X"CB",X"0E",X"7E",X"20",X"1D",X"01",X"F0",
		X"00",X"FD",X"CB",X"0E",X"76",X"28",X"03",X"01",X"80",X"00",X"FD",X"56",X"01",X"1E",X"00",X"CD",
		X"EF",X"55",X"FD",X"74",X"05",X"FD",X"36",X"04",X"C0",X"18",X"25",X"FD",X"7E",X"01",X"FD",X"77",
		X"1B",X"FD",X"36",X"06",X"80",X"FD",X"7E",X"0C",X"FD",X"77",X"18",X"FD",X"36",X"17",X"00",X"67",
		X"2E",X"00",X"FD",X"46",X"01",X"0E",X"00",X"CD",X"10",X"56",X"FD",X"73",X"19",X"FD",X"72",X"1A",
		X"FD",X"7E",X"0F",X"E6",X"3F",X"DD",X"E5",X"E1",X"FD",X"5E",X"10",X"16",X"00",X"19",X"23",X"77",
		X"FD",X"CB",X"0F",X"76",X"28",X"06",X"FD",X"34",X"10",X"C3",X"36",X"54",X"FD",X"36",X"10",X"00",
		X"C9",X"7C",X"F6",X"C4",X"DD",X"77",X"04",X"7D",X"E6",X"0F",X"CD",X"D9",X"55",X"FD",X"77",X"09",
		X"FD",X"36",X"08",X"C0",X"C9",X"FD",X"34",X"1C",X"CD",X"C4",X"55",X"FD",X"7E",X"0E",X"77",X"23",
		X"FD",X"7E",X"0A",X"77",X"23",X"FD",X"7E",X"0B",X"77",X"C9",X"CD",X"C4",X"55",X"35",X"20",X"05",
		X"FD",X"35",X"1C",X"18",X"0A",X"23",X"7E",X"FD",X"77",X"0A",X"23",X"7E",X"FD",X"77",X"0B",X"C9",
		X"FD",X"36",X"02",X"80",X"FD",X"7E",X"0F",X"E6",X"0F",X"07",X"07",X"07",X"FD",X"77",X"11",X"FD",
		X"7E",X"0E",X"E6",X"0F",X"FD",X"77",X"12",X"FD",X"96",X"0C",X"30",X"06",X"FD",X"CB",X"02",X"EE",
		X"ED",X"44",X"67",X"2E",X"00",X"FD",X"46",X"11",X"0E",X"00",X"CD",X"10",X"56",X"FD",X"CB",X"02",
		X"6E",X"28",X"07",X"21",X"00",X"00",X"AF",X"ED",X"52",X"EB",X"FD",X"73",X"15",X"FD",X"72",X"16",
		X"FD",X"7E",X"0C",X"FD",X"77",X"14",X"FD",X"36",X"13",X"00",X"C9",X"FD",X"36",X"00",X"00",X"C9",
		X"FD",X"6E",X"0A",X"FD",X"66",X"0B",X"CF",X"FD",X"73",X"0A",X"FD",X"72",X"0B",X"FD",X"75",X"0E",
		X"FD",X"74",X"0F",X"C9",X"FD",X"E5",X"E1",X"01",X"1D",X"00",X"09",X"FD",X"7E",X"1C",X"87",X"FD",
		X"86",X"1C",X"D6",X"03",X"4F",X"06",X"00",X"09",X"C9",X"3D",X"87",X"5F",X"16",X"00",X"21",X"B7",
		X"52",X"19",X"CF",X"E5",X"C1",X"FD",X"56",X"0D",X"1E",X"00",X"CD",X"EF",X"55",X"7C",X"C9",X"D5",
		X"21",X"00",X"00",X"78",X"A7",X"28",X"0A",X"CB",X"3F",X"30",X"01",X"19",X"EB",X"29",X"EB",X"18",
		X"F3",X"D1",X"79",X"CB",X"3A",X"CB",X"1B",X"A7",X"C8",X"CB",X"27",X"30",X"F6",X"19",X"18",X"F3",
		X"FD",X"E5",X"FD",X"21",X"00",X"00",X"11",X"00",X"01",X"78",X"B1",X"28",X"18",X"AF",X"ED",X"42",
		X"38",X"04",X"FD",X"19",X"18",X"F7",X"09",X"CB",X"38",X"CB",X"19",X"78",X"B1",X"28",X"06",X"CB",
		X"3A",X"CB",X"1B",X"30",X"E8",X"FD",X"E5",X"D1",X"FD",X"E1",X"C9",X"FD",X"35",X"0F",X"20",X"0B",
		X"FD",X"7E",X"10",X"FD",X"77",X"0A",X"FD",X"36",X"00",X"00",X"C9",X"FD",X"6E",X"11",X"FD",X"66",
		X"12",X"FD",X"5E",X"13",X"FD",X"56",X"14",X"19",X"FD",X"75",X"11",X"FD",X"74",X"12",X"7C",X"E6",
		X"0F",X"FD",X"77",X"0A",X"47",X"DD",X"7E",X"00",X"A7",X"28",X"03",X"DD",X"70",X"00",X"FD",X"7E",
		X"0B",X"FD",X"77",X"01",X"FD",X"CB",X"00",X"F6",X"C9",X"DD",X"36",X"00",X"00",X"FD",X"36",X"00",
		X"00",X"C9",X"FD",X"35",X"15",X"20",X"05",X"FD",X"36",X"00",X"00",X"C9",X"FD",X"6E",X"11",X"FD",
		X"66",X"12",X"FD",X"5E",X"13",X"FD",X"56",X"14",X"AF",X"ED",X"52",X"FD",X"75",X"11",X"FD",X"74",
		X"12",X"7C",X"E6",X"0F",X"DD",X"77",X"00",X"A7",X"28",X"DD",X"C9",X"DD",X"36",X"04",X"00",X"FD",
		X"36",X"00",X"00",X"C9",X"DD",X"CB",X"01",X"EE",X"DD",X"6E",X"00",X"26",X"00",X"29",X"11",X"D0",
		X"56",X"19",X"CF",X"4E",X"23",X"06",X"00",X"DD",X"E5",X"D1",X"13",X"13",X"13",X"ED",X"B0",X"C9",
		X"04",X"57",X"1B",X"57",X"32",X"57",X"49",X"57",X"60",X"57",X"69",X"57",X"71",X"57",X"77",X"57",
		X"7D",X"57",X"88",X"57",X"90",X"57",X"9C",X"57",X"B9",X"57",X"B0",X"57",X"A7",X"57",X"C2",X"57",
		X"C8",X"57",X"D7",X"57",X"E0",X"57",X"E8",X"57",X"F7",X"57",X"04",X"58",X"13",X"58",X"00",X"00",
		X"00",X"00",X"1D",X"58",X"16",X"80",X"00",X"00",X"07",X"C0",X"0F",X"AD",X"01",X"00",X"06",X"C0",
		X"0F",X"F0",X"60",X"00",X"60",X"00",X"FF",X"FF",X"01",X"FE",X"18",X"16",X"80",X"00",X"00",X"07",
		X"C0",X"0F",X"00",X"00",X"00",X"07",X"C0",X"0F",X"F0",X"60",X"00",X"60",X"00",X"FD",X"FF",X"01",
		X"FC",X"18",X"16",X"00",X"01",X"00",X"03",X"C0",X"0F",X"AD",X"01",X"00",X"07",X"C0",X"0F",X"F0",
		X"60",X"00",X"60",X"00",X"FD",X"FF",X"01",X"FB",X"08",X"16",X"10",X"00",X"00",X"07",X"C0",X"0F",
		X"AD",X"01",X"00",X"07",X"C0",X"0F",X"C0",X"80",X"00",X"00",X"00",X"FD",X"FF",X"01",X"FD",X"08",
		X"08",X"00",X"00",X"0A",X"07",X"C0",X"0F",X"02",X"BF",X"07",X"01",X"00",X"0F",X"40",X"00",X"0F",
		X"40",X"05",X"00",X"00",X"0F",X"55",X"FA",X"05",X"01",X"00",X"0F",X"55",X"AF",X"0A",X"AD",X"01",
		X"0F",X"60",X"F0",X"59",X"56",X"FA",X"FF",X"FF",X"07",X"04",X"00",X"00",X"07",X"C0",X"0F",X"F0",
		X"0B",X"20",X"00",X"0F",X"9C",X"00",X"0F",X"30",X"00",X"00",X"00",X"00",X"0A",X"00",X"00",X"0F",
		X"60",X"F0",X"50",X"94",X"FE",X"FF",X"FD",X"08",X"04",X"00",X"0A",X"07",X"C0",X"0A",X"DD",X"ED",
		X"08",X"FF",X"00",X"08",X"07",X"C0",X"0B",X"FF",X"1F",X"08",X"7D",X"00",X"0C",X"3E",X"00",X"0C",
		X"38",X"00",X"05",X"E8",X"00",X"0F",X"02",X"7F",X"0E",X"40",X"01",X"0E",X"42",X"01",X"0E",X"0D",
		X"0D",X"40",X"01",X"18",X"41",X"01",X"18",X"08",X"A0",X"03",X"0F",X"E2",X"03",X"0F",X"F0",X"00",
		X"07",X"02",X"00",X"0F",X"06",X"C0",X"0F",X"F0",X"0E",X"D0",X"03",X"0A",X"D1",X"03",X"0A",X"09",
		X"09",X"D0",X"03",X"10",X"D1",X"03",X"10",X"0C",X"98",X"00",X"0F",X"98",X"00",X"0F",X"A0",X"A0",
		X"00",X"38",X"00",X"F0",X"0E",X"20",X"00",X"0A",X"21",X"00",X"0A",X"03",X"01",X"20",X"00",X"10",
		X"21",X"00",X"10",X"09",X"60",X"00",X"0F",X"61",X"00",X"0F",X"60",X"01",X"F0",X"08",X"00",X"00",
		X"00",X"07",X"C0",X"0F",X"01",X"FF",X"DD",X"CB",X"01",X"6E",X"20",X"12",X"CD",X"B4",X"56",X"DD",
		X"7E",X"18",X"DD",X"77",X"02",X"DD",X"CB",X"01",X"F6",X"DD",X"CB",X"01",X"E6",X"C9",X"DD",X"CB",
		X"01",X"66",X"28",X"1D",X"DD",X"6E",X"10",X"DD",X"66",X"11",X"DD",X"75",X"03",X"DD",X"74",X"04",
		X"DD",X"6E",X"12",X"DD",X"66",X"13",X"DD",X"75",X"09",X"DD",X"74",X"0A",X"DD",X"CB",X"01",X"A6",
		X"C9",X"DD",X"7E",X"08",X"A7",X"20",X"04",X"CD",X"9E",X"52",X"C9",X"DD",X"6E",X"03",X"DD",X"66",
		X"04",X"DD",X"5E",X"14",X"DD",X"56",X"15",X"19",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"7E",
		X"16",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",X"0A",X"DD",X"77",X"09",X"DD",X"7E",X"0F",X"DD",
		X"86",X"17",X"DD",X"77",X"0F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"08",
		X"DD",X"77",X"0E",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"09",X"CD",X"B4",X"56",X"21",X"1D",X"6C",
		X"CB",X"D6",X"C9",X"DD",X"7E",X"09",X"DD",X"86",X"03",X"DD",X"A6",X"0A",X"DD",X"77",X"03",X"C0",
		X"CD",X"9E",X"52",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"0A",X"CD",X"B4",X"56",X"21",X"1D",X"6C",
		X"CB",X"D6",X"18",X"2A",X"DD",X"7E",X"09",X"A7",X"20",X"04",X"CD",X"9E",X"52",X"C9",X"DD",X"6E",
		X"03",X"DD",X"66",X"04",X"11",X"09",X"00",X"19",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"6E",
		X"06",X"DD",X"66",X"07",X"19",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"35",X"09",X"DD",X"CB",
		X"01",X"F6",X"DD",X"36",X"02",X"04",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"B4",X"56",
		X"C9",X"DD",X"7E",X"06",X"DD",X"86",X"03",X"DD",X"A6",X"07",X"DD",X"77",X"03",X"C0",X"CD",X"9E",
		X"52",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"B4",X"56",X"C9",X"DD",X"7E",X"06",X"DD",
		X"BE",X"08",X"38",X"12",X"28",X"10",X"DD",X"7E",X"03",X"DD",X"86",X"09",X"30",X"03",X"DD",X"34",
		X"04",X"DD",X"77",X"03",X"18",X"13",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"DD",X"4E",X"0A",X"DD",
		X"46",X"0B",X"09",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"35",X"06",X"DD",X"7E",X"07",X"DD",
		X"86",X"0C",X"DD",X"77",X"07",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"05",
		X"20",X"03",X"CD",X"9E",X"52",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"0C",X"DD",X"CB",X"01",X"F6",
		X"DD",X"36",X"02",X"0B",X"CD",X"B4",X"56",X"C9",X"DD",X"36",X"03",X"0F",X"DD",X"7E",X"08",X"A7",
		X"20",X"04",X"CD",X"9E",X"52",X"C9",X"DD",X"35",X"09",X"DD",X"35",X"09",X"DD",X"7E",X"09",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"08",X"C9",X"DD",X"CB",X"01",X"6E",X"20",
		X"05",X"CD",X"B4",X"56",X"18",X"3B",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"11",X"E0",X"FF",X"19",
		X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"35",X"09",X"20",X"04",X"CD",X"9E",X"52",X"C9",X"DD",
		X"6E",X"06",X"DD",X"66",X"07",X"DD",X"5E",X"0B",X"DD",X"56",X"0C",X"19",X"DD",X"75",X"06",X"DD",
		X"74",X"07",X"DD",X"35",X"0A",X"C0",X"DD",X"7E",X"0D",X"C6",X"03",X"DD",X"77",X"0D",X"FE",X"0C",
		X"D0",X"DD",X"5E",X"0D",X"16",X"00",X"21",X"09",X"5A",X"19",X"7E",X"DD",X"77",X"0A",X"23",X"7E",
		X"DD",X"77",X"0B",X"23",X"7E",X"DD",X"77",X"0C",X"C9",X"05",X"F6",X"FF",X"06",X"06",X"00",X"07",
		X"F0",X"FF",X"FF",X"7C",X"00",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"B4",X"56",X"C9",X"DD",
		X"7E",X"09",X"A7",X"20",X"05",X"DD",X"CB",X"01",X"AE",X"C9",X"DD",X"35",X"09",X"DD",X"7E",X"09",
		X"FE",X"3E",X"38",X"11",X"28",X"0F",X"DD",X"7E",X"03",X"C6",X"1E",X"30",X"03",X"DD",X"34",X"04",
		X"DD",X"77",X"03",X"18",X"10",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"01",X"F9",X"FF",X"09",X"DD",
		X"75",X"03",X"DD",X"74",X"04",X"DD",X"7E",X"0A",X"FE",X"10",X"30",X"0F",X"DD",X"7E",X"06",X"C6",
		X"09",X"30",X"03",X"DD",X"34",X"07",X"DD",X"77",X"06",X"18",X"10",X"DD",X"6E",X"06",X"DD",X"66",
		X"07",X"01",X"FD",X"FF",X"09",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"34",X"0A",X"C9",X"DD",
		X"CB",X"01",X"6E",X"20",X"04",X"CD",X"B4",X"56",X"C9",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"DD",
		X"4E",X"09",X"06",X"00",X"CB",X"79",X"28",X"01",X"05",X"09",X"DD",X"75",X"03",X"DD",X"74",X"04",
		X"DD",X"5E",X"0B",X"DD",X"56",X"0C",X"EB",X"AF",X"ED",X"52",X"F2",X"B4",X"5A",X"11",X"00",X"00",
		X"EB",X"AF",X"ED",X"52",X"DD",X"5E",X"0D",X"16",X"00",X"AF",X"ED",X"52",X"28",X"09",X"FA",X"C7",
		X"5A",X"79",X"ED",X"44",X"DD",X"77",X"09",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"DD",X"4E",X"0A",
		X"06",X"00",X"CB",X"79",X"28",X"01",X"05",X"09",X"DD",X"75",X"06",X"DD",X"74",X"07",X"DD",X"5E",
		X"0E",X"DD",X"56",X"0F",X"EB",X"AF",X"ED",X"52",X"F2",X"F2",X"5A",X"11",X"00",X"00",X"EB",X"AF",
		X"ED",X"52",X"DD",X"5E",X"10",X"16",X"00",X"AF",X"ED",X"52",X"28",X"09",X"FA",X"05",X"5B",X"79",
		X"ED",X"44",X"DD",X"77",X"0A",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"B4",X"56",X"C9",
		X"DD",X"7E",X"0A",X"FE",X"10",X"30",X"1F",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"11",X"FD",X"FF",
		X"19",X"DD",X"75",X"03",X"DD",X"74",X"04",X"DD",X"7E",X"06",X"C6",X"02",X"30",X"03",X"DD",X"34",
		X"07",X"DD",X"77",X"06",X"18",X"1D",X"DD",X"7E",X"03",X"C6",X"02",X"30",X"03",X"DD",X"34",X"04",
		X"DD",X"77",X"03",X"DD",X"6E",X"06",X"DD",X"66",X"07",X"11",X"FE",X"FF",X"19",X"DD",X"75",X"06",
		X"DD",X"74",X"07",X"DD",X"7E",X"09",X"C6",X"FE",X"DD",X"77",X"09",X"CB",X"3F",X"CB",X"3F",X"CB",
		X"3F",X"CB",X"3F",X"DD",X"77",X"05",X"DD",X"77",X"08",X"DD",X"34",X"0A",X"DD",X"7E",X"0A",X"FE",
		X"50",X"38",X"05",X"28",X"03",X"CD",X"9E",X"52",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"0C",X"DD",
		X"CB",X"01",X"F6",X"DD",X"36",X"02",X"0A",X"CD",X"B4",X"56",X"C9",X"DD",X"36",X"03",X"01",X"DD",
		X"7E",X"05",X"A7",X"20",X"04",X"CD",X"9E",X"52",X"C9",X"DD",X"7E",X"09",X"D6",X"08",X"DD",X"77",
		X"09",X"A7",X"1F",X"1F",X"1F",X"1F",X"DD",X"77",X"05",X"DD",X"77",X"08",X"C9",X"DD",X"CB",X"01",
		X"6E",X"20",X"08",X"DD",X"36",X"0F",X"FF",X"CD",X"B4",X"56",X"C9",X"DD",X"7E",X"0F",X"A7",X"20",
		X"04",X"CD",X"9E",X"52",X"C9",X"DD",X"7E",X"09",X"A7",X"20",X"05",X"DD",X"35",X"0F",X"18",X"E7",
		X"DD",X"35",X"09",X"DD",X"7E",X"05",X"A7",X"28",X"14",X"DD",X"35",X"0E",X"DD",X"7E",X"0E",X"CB",
		X"3F",X"CB",X"3F",X"CB",X"3F",X"CB",X"3F",X"DD",X"77",X"05",X"DD",X"77",X"08",X"DD",X"4E",X"0A",
		X"DD",X"46",X"0B",X"DD",X"6E",X"03",X"DD",X"66",X"04",X"09",X"DD",X"75",X"03",X"DD",X"74",X"04",
		X"11",X"20",X"01",X"AF",X"ED",X"52",X"F2",X"10",X"5C",X"EB",X"21",X"00",X"00",X"AF",X"ED",X"52",
		X"11",X"33",X"00",X"AF",X"ED",X"52",X"FA",X"27",X"5C",X"28",X"0C",X"21",X"00",X"00",X"AF",X"ED",
		X"42",X"DD",X"75",X"0A",X"DD",X"74",X"0B",X"DD",X"4E",X"0C",X"DD",X"46",X"0D",X"DD",X"6E",X"06",
		X"DD",X"66",X"07",X"09",X"DD",X"75",X"06",X"DD",X"74",X"07",X"11",X"60",X"00",X"AF",X"ED",X"52",
		X"F2",X"4A",X"5C",X"EB",X"21",X"00",X"00",X"AF",X"ED",X"52",X"11",X"CC",X"0C",X"AF",X"ED",X"52",
		X"FA",X"61",X"5C",X"28",X"0C",X"AF",X"21",X"00",X"00",X"ED",X"42",X"DD",X"75",X"0C",X"DD",X"74",
		X"0D",X"C9",X"DD",X"CB",X"01",X"6E",X"20",X"04",X"CD",X"B4",X"56",X"C9",X"DD",X"7E",X"09",X"DD",
		X"B6",X"0A",X"20",X"02",X"18",X"F2",X"DD",X"7E",X"09",X"D6",X"01",X"30",X"03",X"DD",X"35",X"0A",
		X"DD",X"77",X"09",X"DD",X"7E",X"05",X"A7",X"C8",X"DD",X"35",X"0B",X"DD",X"7E",X"0B",X"A7",X"1F",
		X"1F",X"1F",X"1F",X"DD",X"77",X"05",X"DD",X"77",X"08",X"C9",X"03",X"0F",X"02",X"90",X"00",X"50",
		X"45",X"1C",X"00",X"50",X"03",X"1C",X"00",X"50",X"03",X"1C",X"00",X"50",X"07",X"1C",X"00",X"54",
		X"45",X"20",X"00",X"50",X"03",X"1C",X"00",X"54",X"03",X"20",X"00",X"57",X"07",X"23",X"00",X"A0",
		X"00",X"57",X"45",X"23",X"00",X"58",X"45",X"24",X"00",X"57",X"45",X"23",X"00",X"58",X"45",X"24",
		X"00",X"57",X"45",X"23",X"00",X"58",X"45",X"24",X"00",X"57",X"45",X"23",X"00",X"58",X"45",X"24",
		X"00",X"57",X"45",X"23",X"00",X"57",X"03",X"23",X"00",X"57",X"03",X"23",X"00",X"57",X"45",X"23",
		X"00",X"57",X"45",X"23",X"00",X"57",X"07",X"23",X"07",X"00",X"FF",X"FF",X"00",X"00",X"00",X"00",
		X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"0F",X"02",X"90",X"00",
		X"50",X"87",X"04",X"00",X"50",X"87",X"04",X"00",X"54",X"87",X"08",X"00",X"54",X"87",X"08",X"00",
		X"A0",X"00",X"55",X"87",X"09",X"00",X"55",X"87",X"09",X"00",X"52",X"87",X"07",X"00",X"52",X"87",
		X"07",X"00",X"54",X"87",X"08",X"00",X"54",X"87",X"08",X"00",X"50",X"87",X"04",X"07",X"00",X"FF",
		X"FF",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",X"00",
		X"00",X"05",X"0F",X"02",X"90",X"00",X"5C",X"85",X"23",X"00",X"5C",X"03",X"23",X"00",X"5C",X"03",
		X"23",X"00",X"57",X"85",X"1C",X"00",X"5C",X"85",X"20",X"00",X"A0",X"00",X"5B",X"03",X"20",X"00",
		X"5A",X"03",X"1F",X"00",X"59",X"03",X"1E",X"00",X"58",X"03",X"1D",X"00",X"57",X"03",X"1C",X"00",
		X"58",X"03",X"1D",X"00",X"59",X"03",X"1E",X"00",X"5A",X"03",X"1F",X"00",X"5B",X"45",X"20",X"00",
		X"60",X"45",X"23",X"00",X"5C",X"85",X"17",X"05",X"00",X"FF",X"FF",X"00",X"00",X"0F",X"02",X"90",
		X"85",X"14",X"85",X"16",X"85",X"14",X"85",X"10",X"00",X"A0",X"45",X"10",X"45",X"0F",X"45",X"0D",
		X"45",X"0F",X"87",X"10",X"07",X"00",X"FF",X"FF",X"43",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",
		X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF",X"FF");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
