library ieee;
use ieee.std_logic_1164.all,ieee.numeric_std.all;

entity rom_cpu2 is
port (
	clk  : in  std_logic;
	addr : in  std_logic_vector(12 downto 0);
	data : out std_logic_vector(7 downto 0)
);
end entity;

architecture prom of rom_cpu2 is
	type rom is array(0 to  8191) of std_logic_vector(7 downto 0);
	signal rom_data: rom := (
		X"2A",X"04",X"4B",X"03",X"2C",X"04",X"4D",X"03",X"2E",X"04",X"2E",X"07",X"2D",X"07",X"2C",X"06",
		X"2A",X"02",X"48",X"07",X"29",X"06",X"27",X"00",X"28",X"01",X"49",X"03",X"2A",X"04",X"2B",X"01",
		X"2B",X"00",X"2B",X"06",X"2A",X"06",X"29",X"06",X"28",X"02",X"27",X"00",X"27",X"02",X"00",X"38",
		X"00",X"38",X"12",X"03",X"12",X"04",X"12",X"02",X"13",X"02",X"14",X"05",X"14",X"06",X"15",X"02",
		X"16",X"02",X"17",X"02",X"17",X"01",X"16",X"01",X"15",X"01",X"14",X"01",X"14",X"02",X"15",X"02",
		X"16",X"02",X"17",X"02",X"18",X"00",X"18",X"00",X"17",X"01",X"17",X"00",X"17",X"00",X"14",X"01",
		X"12",X"03",X"12",X"04",X"12",X"02",X"13",X"02",X"14",X"02",X"16",X"02",X"17",X"02",X"18",X"00",
		X"18",X"00",X"17",X"01",X"16",X"01",X"14",X"01",X"13",X"01",X"13",X"05",X"13",X"06",X"15",X"02",
		X"16",X"02",X"18",X"00",X"18",X"00",X"16",X"01",X"15",X"01",X"14",X"01",X"13",X"01",X"12",X"01",
		X"12",X"02",X"13",X"02",X"15",X"02",X"16",X"02",X"16",X"01",X"15",X"03",X"15",X"04",X"16",X"02",
		X"17",X"02",X"00",X"4E",X"00",X"4E",X"17",X"01",X"16",X"01",X"15",X"01",X"14",X"01",X"13",X"01",
		X"12",X"03",X"12",X"04",X"14",X"02",X"15",X"02",X"16",X"02",X"17",X"02",X"18",X"00",X"18",X"00",
		X"17",X"01",X"16",X"01",X"15",X"01",X"13",X"01",X"12",X"01",X"12",X"02",X"13",X"02",X"15",X"02",
		X"16",X"02",X"17",X"02",X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"17",X"00",X"16",X"01",
		X"15",X"01",X"15",X"00",X"14",X"01",X"14",X"00",X"13",X"01",X"13",X"00",X"13",X"02",X"14",X"02",
		X"15",X"02",X"16",X"02",X"17",X"00",X"17",X"02",X"18",X"00",X"17",X"01",X"15",X"01",X"14",X"01",
		X"12",X"03",X"12",X"04",X"12",X"06",X"13",X"00",X"13",X"02",X"12",X"03",X"13",X"02",X"14",X"02",
		X"15",X"00",X"15",X"02",X"16",X"00",X"16",X"00",X"15",X"01",X"14",X"01",X"13",X"01",X"13",X"00",
		X"13",X"02",X"14",X"05",X"14",X"06",X"16",X"00",X"16",X"00",X"15",X"01",X"14",X"01",X"13",X"01",
		X"12",X"03",X"12",X"04",X"12",X"02",X"13",X"02",X"15",X"02",X"16",X"00",X"15",X"01",X"14",X"01",
		X"13",X"01",X"00",X"4E",X"00",X"4E",X"27",X"01",X"27",X"00",X"27",X"00",X"28",X"01",X"28",X"00",
		X"49",X"03",X"2A",X"04",X"2B",X"01",X"2B",X"00",X"2C",X"03",X"2C",X"02",X"4A",X"07",X"2B",X"06",
		X"2A",X"03",X"49",X"07",X"2A",X"06",X"28",X"07",X"27",X"00",X"28",X"01",X"29",X"01",X"29",X"07",
		X"28",X"07",X"27",X"00",X"27",X"00",X"28",X"01",X"28",X"07",X"27",X"00",X"27",X"00",X"28",X"01",
		X"29",X"04",X"2A",X"03",X"2B",X"01",X"2C",X"03",X"2D",X"01",X"2D",X"07",X"2C",X"07",X"2B",X"07",
		X"2A",X"02",X"29",X"02",X"28",X"02",X"28",X"00",X"27",X"02",X"20",X"27",X"01",X"27",X"00",X"27",
		X"00",X"27",X"00",X"28",X"01",X"28",X"00",X"29",X"01",X"2A",X"01",X"4B",X"03",X"2C",X"04",X"2C",
		X"00",X"2C",X"07",X"2B",X"07",X"2A",X"07",X"29",X"00",X"29",X"02",X"27",X"00",X"27",X"00",X"27",
		X"00",X"27",X"00",X"27",X"00",X"27",X"00",X"28",X"01",X"29",X"04",X"29",X"07",X"28",X"02",X"27",
		X"00",X"27",X"00",X"28",X"04",X"29",X"09",X"28",X"00",X"28",X"02",X"27",X"02",X"27",X"04",X"28",
		X"01",X"49",X"03",X"2A",X"04",X"2B",X"01",X"2C",X"09",X"2B",X"06",X"00",X"08",X"00",X"08",X"11",
		X"01",X"10",X"01",X"10",X"00",X"11",X"02",X"12",X"02",X"14",X"02",X"16",X"02",X"17",X"02",X"00",
		X"08",X"00",X"08",X"2A",X"02",X"29",X"02",X"28",X"02",X"27",X"00",X"28",X"01",X"29",X"03",X"4A",
		X"03",X"2B",X"04",X"2C",X"04",X"00",X"11",X"00",X"11",X"00",X"08",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"17",X"00",X"15",X"01",X"13",X"01",X"11",X"01",X"0F",X"01",X"0F",X"00",X"0F",
		X"02",X"10",X"02",X"12",X"02",X"13",X"02",X"15",X"02",X"16",X"02",X"17",X"02",X"00",X"11",X"00",
		X"11",X"00",X"03",X"4D",X"03",X"4E",X"05",X"4F",X"05",X"30",X"04",X"31",X"09",X"30",X"07",X"4D",
		X"07",X"4E",X"08",X"2F",X"06",X"2C",X"07",X"2B",X"02",X"2A",X"02",X"29",X"02",X"28",X"00",X"29",
		X"01",X"29",X"00",X"48",X"07",X"29",X"06",X"27",X"00",X"27",X"00",X"27",X"02",X"20",X"20",X"01",
		X"40",X"01",X"40",X"18",X"00",X"17",X"01",X"15",X"01",X"14",X"01",X"13",X"01",X"13",X"00",X"13",
		X"02",X"14",X"02",X"15",X"02",X"16",X"02",X"17",X"02",X"AE",X"17",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"AF",X"17",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"14",X"01",X"13",X"01",X"13",
		X"00",X"13",X"00",X"13",X"02",X"14",X"02",X"15",X"01",X"14",X"01",X"14",X"00",X"14",X"00",X"AF",
		X"15",X"14",X"02",X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"00",X"16",X"02",X"17",X"02",X"18",
		X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"AD",X"17",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"17",X"01",X"17",X"00",X"16",X"01",X"15",X"01",X"14",X"01",X"12",X"01",X"11",
		X"01",X"11",X"00",X"11",X"00",X"11",X"02",X"12",X"02",X"15",X"02",X"16",X"02",X"17",X"00",X"17",
		X"00",X"16",X"01",X"15",X"01",X"AD",X"13",X"14",X"01",X"14",X"00",X"14",X"00",X"14",X"00",X"14",
		X"00",X"13",X"01",X"12",X"01",X"12",X"00",X"12",X"02",X"14",X"02",X"16",X"02",X"18",X"00",X"18",
		X"00",X"18",X"00",X"15",X"01",X"13",X"01",X"12",X"01",X"10",X"01",X"0E",X"01",X"0D",X"00",X"0D",
		X"00",X"0D",X"02",X"0F",X"02",X"11",X"02",X"14",X"02",X"15",X"02",X"17",X"02",X"18",X"00",X"17",
		X"01",X"17",X"00",X"16",X"01",X"15",X"01",X"15",X"00",X"14",X"01",X"13",X"01",X"13",X"00",X"13",
		X"00",X"12",X"01",X"12",X"00",X"11",X"01",X"11",X"00",X"10",X"01",X"10",X"00",X"10",X"00",X"11",
		X"02",X"14",X"02",X"16",X"02",X"17",X"02",X"AE",X"15",X"18",X"00",X"16",X"00",X"16",X"00",X"16",
		X"00",X"15",X"01",X"14",X"01",X"14",X"00",X"AC",X"12",X"13",X"01",X"13",X"00",X"13",X"00",X"13",
		X"00",X"13",X"02",X"14",X"00",X"14",X"02",X"15",X"02",X"17",X"02",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"14",X"01",X"13",X"01",X"11",X"01",X"10",X"01",X"10",
		X"00",X"10",X"00",X"10",X"02",X"13",X"02",X"16",X"02",X"17",X"02",X"17",X"01",X"16",X"01",X"AE",
		X"14",X"15",X"01",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"00",X"14",X"01",X"13",X"01",X"12",
		X"01",X"12",X"00",X"12",X"02",X"15",X"02",X"16",X"02",X"AD",X"17",X"17",X"02",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"16",X"00",X"16",X"00",X"AE",X"14",X"15",
		X"01",X"15",X"00",X"15",X"00",X"15",X"00",X"15",X"02",X"18",X"00",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"16",X"01",X"15",X"01",X"15",X"00",X"15",
		X"00",X"15",X"02",X"AE",X"17",X"16",X"02",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"17",
		X"01",X"16",X"01",X"16",X"00",X"15",X"01",X"14",X"01",X"14",X"00",X"14",X"00",X"13",X"01",X"12",
		X"01",X"12",X"00",X"11",X"01",X"10",X"01",X"10",X"00",X"0F",X"01",X"0F",X"00",X"11",X"02",X"12",
		X"02",X"15",X"02",X"16",X"02",X"17",X"02",X"18",X"00",X"AE",X"17",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"14",X"01",X"14",X"00",X"16",
		X"02",X"17",X"00",X"AF",X"16",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"00",X"17",X"02",X"17",
		X"01",X"16",X"01",X"14",X"01",X"14",X"00",X"14",X"00",X"14",X"02",X"17",X"02",X"18",X"00",X"AD",
		X"17",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"14",
		X"01",X"14",X"00",X"13",X"01",X"13",X"00",X"13",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"AE",X"16",X"17",X"00",X"17",X"00",X"17",
		X"00",X"17",X"00",X"16",X"01",X"15",X"01",X"13",X"01",X"13",X"00",X"13",X"00",X"18",X"00",X"18",
		X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"14",X"01",X"13",X"01",X"10",X"01",X"0E",X"01",X"0D",
		X"01",X"0D",X"00",X"0D",X"02",X"0E",X"02",X"10",X"02",X"15",X"02",X"16",X"02",X"18",X"00",X"18",
		X"00",X"17",X"01",X"15",X"01",X"14",X"01",X"14",X"00",X"14",X"02",X"16",X"02",X"16",X"01",X"AC",
		X"13",X"14",X"01",X"14",X"00",X"14",X"00",X"14",X"00",X"14",X"02",X"15",X"00",X"15",X"00",X"13",
		X"01",X"12",X"01",X"12",X"00",X"12",X"00",X"12",X"02",X"14",X"02",X"15",X"02",X"AD",X"17",X"17",
		X"02",X"18",X"00",X"18",X"00",X"18",X"00",X"18",X"00",X"17",X"01",X"16",X"01",X"15",X"01",X"15",
		X"00",X"15",X"02",X"17",X"02",X"00",X"20",X"00",X"20",X"18",X"01",X"17",X"01",X"16",X"01",X"15",
		X"01",X"14",X"01",X"13",X"01",X"12",X"01",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",
		X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",
		X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"00",X"12",X"02",X"13",X"02",X"14",
		X"02",X"15",X"02",X"16",X"02",X"17",X"02",X"18",X"02",X"00",X"20",X"00",X"20",X"27",X"03",X"28",
		X"03",X"29",X"03",X"2A",X"03",X"2B",X"03",X"2C",X"03",X"2D",X"03",X"2D",X"00",X"2D",X"00",X"2D",
		X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",
		X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",X"00",X"2D",
		X"04",X"2C",X"04",X"2B",X"04",X"2A",X"04",X"29",X"04",X"28",X"04",X"27",X"04",X"A5",X"25",X"D5",
		X"25",X"07",X"26",X"31",X"26",X"00",X"60",X"40",X"A0",X"41",X"A1",X"42",X"62",X"03",X"23",X"40",
		X"A4",X"41",X"A5",X"42",X"66",X"43",X"27",X"64",X"28",X"40",X"A9",X"41",X"AA",X"42",X"6B",X"43",
		X"2C",X"64",X"2D",X"40",X"AE",X"41",X"AF",X"42",X"70",X"43",X"31",X"64",X"32",X"40",X"B3",X"41",
		X"B4",X"42",X"75",X"83",X"36",X"00",X"CD",X"41",X"20",X"42",X"41",X"03",X"42",X"40",X"23",X"41",
		X"24",X"42",X"45",X"43",X"46",X"44",X"27",X"65",X"28",X"40",X"29",X"41",X"2A",X"42",X"4B",X"43",
		X"4C",X"44",X"2D",X"65",X"2E",X"40",X"2F",X"41",X"30",X"42",X"51",X"43",X"52",X"44",X"33",X"65",
		X"34",X"41",X"35",X"42",X"56",X"83",X"57",X"00",X"87",X"40",X"A0",X"41",X"A1",X"42",X"A2",X"43",
		X"63",X"04",X"24",X"40",X"A5",X"41",X"A6",X"42",X"A7",X"43",X"68",X"04",X"29",X"40",X"AA",X"41",
		X"AB",X"42",X"AC",X"43",X"6D",X"04",X"2E",X"40",X"AF",X"41",X"B0",X"42",X"B1",X"43",X"72",X"84",
		X"33",X"00",X"B3",X"41",X"A0",X"02",X"C1",X"40",X"A2",X"41",X"A3",X"42",X"C4",X"43",X"C5",X"64",
		X"86",X"40",X"A7",X"41",X"A8",X"42",X"C9",X"43",X"CA",X"64",X"8B",X"40",X"AC",X"41",X"AD",X"42",
		X"CE",X"43",X"CF",X"64",X"90",X"41",X"B1",X"82",X"D2",X"DD",X"CB",X"00",X"66",X"C2",X"50",X"28",
		X"DD",X"CB",X"00",X"6E",X"20",X"3B",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"02",X"00",X"DD",X"36",
		X"03",X"38",X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"40",X"DD",X"36",X"06",X"00",X"DD",X"36",
		X"07",X"00",X"DD",X"36",X"08",X"00",X"DD",X"36",X"09",X"00",X"DD",X"36",X"0A",X"00",X"DD",X"36",
		X"0B",X"00",X"DD",X"36",X"01",X"40",X"3A",X"1D",X"6C",X"A7",X"C0",X"1E",X"19",X"CD",X"FB",X"06",
		X"C9",X"DD",X"CB",X"00",X"4E",X"20",X"2B",X"FD",X"7E",X"1E",X"47",X"FD",X"AE",X"28",X"E6",X"60",
		X"C0",X"CB",X"70",X"28",X"08",X"DD",X"CB",X"00",X"C6",X"DD",X"36",X"05",X"80",X"DD",X"CB",X"00",
		X"CE",X"FD",X"35",X"00",X"CD",X"AF",X"09",X"2A",X"DD",X"60",X"22",X"7C",X"60",X"21",X"00",X"60",
		X"CB",X"F6",X"DD",X"CB",X"00",X"5E",X"20",X"1C",X"3A",X"1D",X"6C",X"A7",X"20",X"16",X"DD",X"CB",
		X"00",X"DE",X"DD",X"CB",X"00",X"46",X"20",X"07",X"1E",X"13",X"CD",X"FB",X"06",X"18",X"05",X"1E",
		X"16",X"CD",X"FB",X"06",X"CD",X"51",X"29",X"2F",X"E6",X"05",X"28",X"37",X"CB",X"57",X"20",X"05",
		X"11",X"80",X"FE",X"18",X"03",X"11",X"80",X"01",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"19",X"7C",
		X"FE",X"78",X"30",X"1F",X"FE",X"38",X"38",X"1B",X"DD",X"74",X"03",X"DD",X"75",X"04",X"7C",X"D6",
		X"38",X"57",X"ED",X"4B",X"DF",X"60",X"CD",X"3C",X"3A",X"ED",X"5B",X"DD",X"60",X"19",X"22",X"7C",
		X"60",X"18",X"00",X"CD",X"71",X"29",X"2F",X"E6",X"0A",X"28",X"22",X"CB",X"5F",X"20",X"05",X"21",
		X"00",X"01",X"18",X"03",X"21",X"00",X"FF",X"DD",X"56",X"05",X"DD",X"5E",X"06",X"19",X"7C",X"FE",
		X"C0",X"30",X"0A",X"FE",X"40",X"38",X"06",X"DD",X"74",X"05",X"DD",X"75",X"06",X"3A",X"60",X"63",
		X"17",X"38",X"1F",X"CD",X"98",X"29",X"CB",X"67",X"20",X"18",X"21",X"60",X"63",X"CB",X"FE",X"23",
		X"23",X"EB",X"21",X"56",X"63",X"01",X"05",X"00",X"ED",X"B0",X"EB",X"36",X"00",X"1E",X"04",X"CD",
		X"FB",X"06",X"DD",X"7E",X"0A",X"A7",X"20",X"39",X"21",X"68",X"63",X"CB",X"7E",X"28",X"07",X"21",
		X"79",X"63",X"CB",X"7E",X"20",X"2E",X"EB",X"CD",X"A9",X"29",X"1F",X"38",X"27",X"EB",X"CB",X"FE",
		X"23",X"23",X"EB",X"21",X"56",X"63",X"01",X"05",X"00",X"ED",X"B0",X"EB",X"36",X"00",X"ED",X"5B",
		X"7C",X"60",X"23",X"72",X"23",X"73",X"DD",X"36",X"0A",X"20",X"1E",X"05",X"CD",X"FB",X"06",X"18",
		X"03",X"DD",X"35",X"0A",X"3A",X"03",X"60",X"2F",X"E6",X"03",X"20",X"75",X"06",X"07",X"0E",X"03",
		X"CD",X"60",X"0A",X"28",X"05",X"DD",X"CB",X"00",X"E6",X"C9",X"FD",X"7E",X"1E",X"FD",X"AE",X"28",
		X"E6",X"60",X"28",X"5D",X"DD",X"7E",X"05",X"E6",X"F8",X"5F",X"CD",X"F6",X"0A",X"DD",X"86",X"03",
		X"E6",X"F8",X"57",X"CD",X"03",X"0B",X"11",X"00",X"04",X"DD",X"CB",X"00",X"46",X"20",X"22",X"7E",
		X"FE",X"FF",X"20",X"3D",X"19",X"7E",X"E6",X"07",X"FE",X"06",X"20",X"35",X"DD",X"CB",X"00",X"C6",
		X"1E",X"13",X"CD",X"0E",X"07",X"1E",X"08",X"CD",X"FB",X"06",X"1E",X"16",X"CD",X"FB",X"06",X"18",
		X"20",X"7E",X"FE",X"FF",X"20",X"08",X"19",X"7E",X"E6",X"07",X"FE",X"06",X"28",X"13",X"DD",X"CB",
		X"00",X"86",X"1E",X"16",X"CD",X"0E",X"07",X"1E",X"03",X"CD",X"FB",X"06",X"1E",X"13",X"CD",X"FB",
		X"06",X"06",X"C0",X"0E",X"00",X"16",X"03",X"CD",X"02",X"06",X"06",X"0D",X"CD",X"7A",X"06",X"C9",
		X"CD",X"7B",X"0B",X"DA",X"39",X"29",X"DD",X"7E",X"09",X"FE",X"10",X"D2",X"39",X"29",X"DD",X"34",
		X"09",X"E6",X"0C",X"28",X"0B",X"FE",X"04",X"28",X"25",X"FE",X"08",X"28",X"5A",X"C3",X"00",X"29",
		X"01",X"74",X"C0",X"16",X"03",X"CD",X"02",X"06",X"DD",X"7E",X"09",X"FE",X"01",X"C0",X"1E",X"13",
		X"CD",X"0E",X"07",X"1E",X"16",X"CD",X"0E",X"07",X"1E",X"00",X"CD",X"FB",X"06",X"C9",X"11",X"F8",
		X"F8",X"CD",X"EF",X"0B",X"01",X"78",X"C0",X"16",X"0C",X"CD",X"08",X"06",X"11",X"F8",X"08",X"CD",
		X"EF",X"0B",X"01",X"7C",X"C0",X"16",X"0C",X"CD",X"08",X"06",X"11",X"08",X"F8",X"CD",X"EF",X"0B",
		X"01",X"80",X"C0",X"16",X"0C",X"CD",X"08",X"06",X"11",X"08",X"08",X"CD",X"EF",X"0B",X"01",X"84",
		X"C0",X"16",X"0C",X"CD",X"08",X"06",X"C9",X"11",X"F8",X"F8",X"CD",X"EF",X"0B",X"01",X"88",X"C0",
		X"16",X"02",X"CD",X"08",X"06",X"11",X"F8",X"08",X"CD",X"EF",X"0B",X"01",X"8C",X"C0",X"16",X"02",
		X"CD",X"08",X"06",X"11",X"08",X"F8",X"CD",X"EF",X"0B",X"01",X"8C",X"F0",X"16",X"02",X"CD",X"08",
		X"06",X"11",X"08",X"08",X"CD",X"EF",X"0B",X"01",X"88",X"F0",X"16",X"02",X"CD",X"08",X"06",X"C9",
		X"11",X"F8",X"F8",X"CD",X"EF",X"0B",X"01",X"90",X"C0",X"16",X"0E",X"CD",X"08",X"06",X"11",X"F8",
		X"08",X"CD",X"EF",X"0B",X"01",X"94",X"C0",X"16",X"0E",X"CD",X"08",X"06",X"11",X"08",X"F8",X"CD",
		X"EF",X"0B",X"01",X"94",X"F0",X"16",X"0E",X"CD",X"08",X"06",X"11",X"08",X"08",X"CD",X"EF",X"0B",
		X"01",X"90",X"F0",X"16",X"0E",X"CD",X"08",X"06",X"C9",X"DD",X"36",X"00",X"00",X"21",X"49",X"63",
		X"CB",X"FE",X"21",X"00",X"60",X"CB",X"B6",X"23",X"CB",X"FE",X"21",X"00",X"00",X"22",X"7C",X"60",
		X"C9",X"21",X"00",X"60",X"CB",X"7E",X"28",X"0A",X"3A",X"00",X"90",X"CB",X"46",X"C8",X"3A",X"01",
		X"90",X"C9",X"DD",X"34",X"0B",X"DD",X"CB",X"0B",X"6E",X"20",X"03",X"3E",X"FB",X"C9",X"3E",X"FE",
		X"C9",X"21",X"00",X"60",X"CB",X"7E",X"28",X"0A",X"3A",X"00",X"90",X"CB",X"46",X"C8",X"3A",X"01",
		X"90",X"C9",X"3A",X"A1",X"60",X"DD",X"86",X"03",X"CD",X"EF",X"2B",X"D6",X"30",X"DD",X"BE",X"05",
		X"30",X"03",X"3E",X"F7",X"C9",X"3E",X"FD",X"C9",X"21",X"00",X"60",X"AF",X"CB",X"7E",X"C8",X"3A",
		X"00",X"90",X"CB",X"46",X"C8",X"3A",X"01",X"90",X"C9",X"21",X"00",X"60",X"AF",X"CB",X"7E",X"C8",
		X"3A",X"00",X"E0",X"CB",X"46",X"C8",X"1F",X"C9",X"DD",X"CB",X"00",X"66",X"20",X"4C",X"21",X"00",
		X"08",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"19",X"7C",X"FE",X"F0",X"30",X"61",X"DD",X"74",X"03",
		X"DD",X"75",X"04",X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",X"26",X"0C",X"06",X"18",X"0E",X"09",
		X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",X"0A",X"38",X"17",X"FD",X"19",X"10",X"F2",X"06",X"10",
		X"0E",X"01",X"CD",X"60",X"0A",X"20",X"0E",X"06",X"80",X"0E",X"6C",X"16",X"03",X"CD",X"02",X"06",
		X"C9",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"7E",X"07",X"FE",X"0C",X"30",
		X"1D",X"CD",X"7B",X"0B",X"38",X"18",X"DD",X"7E",X"07",X"21",X"A3",X"0B",X"CD",X"93",X"0B",X"DD",
		X"34",X"07",X"DD",X"7E",X"07",X"FE",X"01",X"C0",X"1E",X"12",X"CD",X"FB",X"06",X"C9",X"DD",X"36",
		X"00",X"00",X"21",X"01",X"60",X"CB",X"FE",X"C9",X"DD",X"CB",X"00",X"66",X"C2",X"C6",X"2B",X"DD",
		X"CB",X"00",X"46",X"C2",X"DA",X"2A",X"21",X"80",X"01",X"DD",X"56",X"05",X"DD",X"5E",X"06",X"19",
		X"DD",X"74",X"05",X"DD",X"75",X"06",X"ED",X"5B",X"7C",X"60",X"DD",X"66",X"08",X"DD",X"6E",X"09",
		X"A7",X"ED",X"52",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"19",X"7C",X"FE",X"08",X"DA",X"B7",X"2B",
		X"FE",X"F8",X"D2",X"B7",X"2B",X"DD",X"74",X"03",X"DD",X"75",X"04",X"06",X"03",X"0E",X"01",X"CD",
		X"60",X"0A",X"28",X"4C",X"3A",X"A1",X"60",X"DD",X"86",X"03",X"CD",X"EF",X"2B",X"D6",X"10",X"DD",
		X"BE",X"05",X"38",X"05",X"DD",X"CB",X"00",X"E6",X"C9",X"DD",X"CB",X"00",X"C6",X"DD",X"36",X"08",
		X"1E",X"C6",X"14",X"DD",X"77",X"0B",X"DD",X"36",X"0C",X"00",X"DD",X"77",X"0F",X"DD",X"36",X"10",
		X"00",X"DD",X"7E",X"03",X"DD",X"77",X"09",X"DD",X"77",X"0D",X"DD",X"7E",X"04",X"DD",X"77",X"0A",
		X"DD",X"77",X"0E",X"1E",X"05",X"CD",X"0E",X"07",X"1E",X"12",X"CD",X"FB",X"06",X"C3",X"A1",X"2B",
		X"06",X"80",X"0E",X"6D",X"16",X"0D",X"CD",X"02",X"06",X"C9",X"DD",X"35",X"08",X"CA",X"BC",X"2B",
		X"3A",X"03",X"60",X"E6",X"03",X"FE",X"01",X"20",X"5C",X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",
		X"06",X"0C",X"CD",X"15",X"0A",X"28",X"23",X"FD",X"7E",X"02",X"A7",X"20",X"1D",X"FD",X"7E",X"00",
		X"E6",X"07",X"FE",X"05",X"28",X"14",X"DD",X"7E",X"09",X"D6",X"0B",X"FD",X"BE",X"03",X"30",X"0A",
		X"DD",X"7E",X"0D",X"C6",X"0B",X"FD",X"BE",X"03",X"30",X"27",X"FD",X"19",X"10",X"D4",X"FD",X"21",
		X"D0",X"64",X"CD",X"15",X"0A",X"28",X"1E",X"FD",X"7E",X"02",X"A7",X"20",X"18",X"DD",X"7E",X"09",
		X"D6",X"0A",X"FD",X"BE",X"03",X"30",X"0E",X"DD",X"7E",X"0D",X"C6",X"0A",X"FD",X"BE",X"03",X"38",
		X"04",X"FD",X"CB",X"00",X"E6",X"ED",X"5B",X"7C",X"60",X"DD",X"7E",X"09",X"FE",X"10",X"38",X"0D",
		X"67",X"DD",X"6E",X"0A",X"A7",X"ED",X"52",X"DD",X"74",X"09",X"DD",X"75",X"0A",X"DD",X"7E",X"0D",
		X"FE",X"10",X"38",X"58",X"67",X"DD",X"6E",X"0E",X"CB",X"2A",X"CB",X"1B",X"A7",X"ED",X"52",X"DD",
		X"74",X"0D",X"DD",X"75",X"0E",X"3A",X"A1",X"60",X"84",X"CD",X"EF",X"2B",X"C6",X"04",X"47",X"DD",
		X"96",X"0F",X"30",X"02",X"ED",X"44",X"FE",X"20",X"30",X"32",X"DD",X"70",X"0F",X"DD",X"CB",X"08",
		X"46",X"20",X"0E",X"DD",X"7E",X"09",X"DD",X"77",X"03",X"DD",X"7E",X"0B",X"DD",X"77",X"05",X"18",
		X"0C",X"DD",X"7E",X"0D",X"DD",X"77",X"03",X"DD",X"7E",X"0F",X"DD",X"77",X"05",X"06",X"C0",X"0E",
		X"BC",X"16",X"05",X"CD",X"02",X"06",X"C9",X"1E",X"05",X"CD",X"0E",X"07",X"DD",X"36",X"00",X"00",
		X"21",X"01",X"60",X"CB",X"FE",X"C9",X"DD",X"7E",X"07",X"A7",X"20",X"0A",X"1E",X"05",X"CD",X"0E",
		X"07",X"1E",X"12",X"CD",X"FB",X"06",X"DD",X"7E",X"07",X"FE",X"0C",X"30",X"DF",X"CD",X"7B",X"0B",
		X"38",X"DA",X"DD",X"7E",X"07",X"21",X"A3",X"0B",X"CD",X"93",X"0B",X"DD",X"34",X"07",X"C9",X"E6",
		X"F8",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"A2",X"60",X"19",X"7E",X"87",X"87",X"87",X"C9",
		X"3A",X"54",X"63",X"17",X"38",X"05",X"DD",X"36",X"00",X"00",X"C9",X"2A",X"78",X"60",X"CD",X"1E",
		X"2C",X"22",X"78",X"60",X"2A",X"7A",X"60",X"CD",X"1E",X"2C",X"22",X"7A",X"60",X"C9",X"11",X"80",
		X"FF",X"19",X"7C",X"FE",X"FD",X"D0",X"FE",X"04",X"D8",X"26",X"03",X"C9",X"DD",X"CB",X"00",X"6E",
		X"20",X"08",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"02",X"0E",X"DD",X"CB",X"02",X"46",X"20",X"19",
		X"DD",X"7E",X"00",X"E6",X"07",X"87",X"5F",X"16",X"00",X"21",X"73",X"2C",X"19",X"5E",X"23",X"56",
		X"EB",X"CD",X"75",X"09",X"CD",X"75",X"09",X"18",X"09",X"21",X"B7",X"D0",X"01",X"02",X"08",X"CD",
		X"82",X"09",X"DD",X"36",X"01",X"08",X"DD",X"35",X"02",X"C0",X"DD",X"36",X"01",X"00",X"DD",X"36",
		X"00",X"00",X"C9",X"81",X"2C",X"90",X"2C",X"A3",X"2C",X"B4",X"2C",X"CA",X"2C",X"DF",X"2C",X"F2",
		X"2C",X"B7",X"D0",X"03",X"1E",X"0F",X"18",X"D9",X"D0",X"06",X"0C",X"18",X"16",X"12",X"17",X"10",
		X"B7",X"D0",X"06",X"11",X"18",X"16",X"12",X"17",X"10",X"D8",X"D0",X"07",X"16",X"12",X"1C",X"1C",
		X"12",X"15",X"0E",X"B7",X"D0",X"05",X"1B",X"0A",X"0D",X"0A",X"1B",X"D9",X"D0",X"06",X"1C",X"0E",
		X"0A",X"1B",X"0C",X"11",X"B7",X"D0",X"08",X"1D",X"11",X"0E",X"24",X"1D",X"0A",X"17",X"14",X"D7",
		X"D0",X"08",X"12",X"1C",X"24",X"0F",X"18",X"1E",X"17",X"0D",X"B7",X"D0",X"07",X"1D",X"11",X"0E",
		X"24",X"1C",X"0E",X"0A",X"D7",X"D0",X"08",X"12",X"1C",X"24",X"0F",X"18",X"1E",X"17",X"0D",X"B7",
		X"D0",X"07",X"16",X"12",X"1C",X"1C",X"12",X"15",X"0E",X"D9",X"D0",X"06",X"0C",X"18",X"16",X"12",
		X"17",X"10",X"B7",X"D0",X"04",X"1C",X"1E",X"0B",X"2D",X"D9",X"D0",X"06",X"16",X"0A",X"1B",X"12",
		X"17",X"0E",X"4E",X"21",X"00",X"60",X"CB",X"76",X"20",X"2B",X"21",X"54",X"63",X"CB",X"7E",X"20",
		X"05",X"DD",X"36",X"00",X"00",X"C9",X"DD",X"CB",X"00",X"6E",X"20",X"19",X"DD",X"CB",X"00",X"EE",
		X"DD",X"36",X"02",X"00",X"DD",X"36",X"04",X"10",X"DD",X"36",X"05",X"00",X"DD",X"36",X"08",X"00",
		X"DD",X"36",X"0A",X"00",X"C9",X"26",X"00",X"DD",X"6E",X"02",X"DD",X"34",X"02",X"DD",X"7E",X"02",
		X"FE",X"07",X"38",X"04",X"DD",X"36",X"02",X"00",X"29",X"11",X"52",X"2D",X"19",X"5E",X"23",X"56",
		X"EB",X"E9",X"60",X"2D",X"03",X"31",X"87",X"32",X"51",X"33",X"A1",X"33",X"1E",X"34",X"B1",X"34",
		X"FD",X"CB",X"2E",X"7E",X"28",X"48",X"CD",X"D8",X"2D",X"7E",X"FE",X"FF",X"28",X"0B",X"CD",X"1E",
		X"2E",X"CD",X"40",X"2E",X"FD",X"34",X"6A",X"18",X"ED",X"FD",X"CB",X"69",X"7E",X"28",X"13",X"CD",
		X"F2",X"2D",X"7E",X"FE",X"FF",X"28",X"0B",X"CD",X"1E",X"2E",X"CD",X"40",X"2E",X"FD",X"34",X"6C",
		X"18",X"ED",X"FD",X"CB",X"2E",X"BE",X"FD",X"7E",X"32",X"FD",X"77",X"69",X"FD",X"36",X"6A",X"00",
		X"CB",X"7F",X"28",X"0A",X"FD",X"7E",X"33",X"FD",X"77",X"6B",X"FD",X"36",X"6C",X"00",X"CD",X"D8",
		X"2D",X"7E",X"FE",X"FF",X"28",X"0B",X"CD",X"0C",X"2E",X"38",X"06",X"CD",X"40",X"2E",X"FD",X"34",
		X"6A",X"FD",X"CB",X"69",X"7E",X"C8",X"CD",X"F2",X"2D",X"7E",X"FE",X"FF",X"C8",X"CD",X"0C",X"2E",
		X"D8",X"CD",X"40",X"2E",X"FD",X"34",X"6C",X"C9",X"FD",X"7E",X"69",X"E6",X"1F",X"87",X"5F",X"16",
		X"00",X"21",X"01",X"2F",X"19",X"5E",X"23",X"56",X"FD",X"7E",X"6A",X"87",X"87",X"6F",X"26",X"00",
		X"19",X"C9",X"FD",X"7E",X"6B",X"E6",X"1F",X"87",X"5F",X"16",X"00",X"21",X"01",X"2F",X"19",X"5E",
		X"23",X"56",X"FD",X"7E",X"6C",X"87",X"87",X"6F",X"26",X"00",X"19",X"C9",X"E5",X"23",X"56",X"23",
		X"5E",X"EB",X"FD",X"56",X"34",X"FD",X"5E",X"35",X"A7",X"ED",X"52",X"EB",X"E1",X"C9",X"CD",X"0C",
		X"2E",X"E5",X"D5",X"FD",X"7E",X"32",X"E6",X"1F",X"87",X"5F",X"16",X"00",X"21",X"82",X"1B",X"19",
		X"5E",X"23",X"56",X"EB",X"56",X"23",X"5E",X"EB",X"29",X"29",X"29",X"D1",X"19",X"EB",X"E1",X"C9",
		X"FD",X"CB",X"69",X"6E",X"C0",X"FD",X"CB",X"69",X"76",X"20",X"05",X"CB",X"66",X"C8",X"18",X"03",
		X"CB",X"5E",X"C8",X"7E",X"E6",X"07",X"FE",X"04",X"20",X"0A",X"D5",X"E5",X"CD",X"75",X"07",X"E1",
		X"D1",X"E6",X"01",X"C8",X"DD",X"E5",X"D5",X"FD",X"E5",X"DD",X"E1",X"11",X"6F",X"00",X"DD",X"19",
		X"11",X"08",X"00",X"06",X"18",X"DD",X"CB",X"00",X"7E",X"28",X"08",X"DD",X"19",X"10",X"F6",X"D1",
		X"DD",X"E1",X"C9",X"D1",X"7E",X"E6",X"07",X"F6",X"80",X"DD",X"77",X"00",X"E5",X"21",X"00",X"04",
		X"A7",X"ED",X"52",X"E5",X"2A",X"8C",X"63",X"55",X"5C",X"2A",X"A0",X"60",X"A7",X"ED",X"52",X"EB",
		X"E1",X"7C",X"65",X"FD",X"6E",X"36",X"A7",X"ED",X"52",X"DE",X"00",X"DD",X"77",X"01",X"DD",X"74",
		X"02",X"DD",X"75",X"03",X"E1",X"23",X"23",X"23",X"FD",X"7E",X"37",X"87",X"87",X"87",X"86",X"DD",
		X"77",X"04",X"DD",X"36",X"05",X"00",X"2A",X"A0",X"60",X"DD",X"74",X"06",X"DD",X"75",X"07",X"DD",
		X"E5",X"E1",X"DD",X"E1",X"7E",X"E6",X"07",X"FE",X"04",X"C8",X"DD",X"7E",X"09",X"A7",X"28",X"04",
		X"DD",X"35",X"09",X"C9",X"CB",X"DE",X"FD",X"7E",X"0B",X"E6",X"30",X"0F",X"0F",X"0F",X"5F",X"16",
		X"00",X"21",X"FB",X"30",X"3A",X"DC",X"60",X"A7",X"28",X"01",X"23",X"19",X"7E",X"DD",X"77",X"09",
		X"C9",X"27",X"2F",X"FA",X"30",X"FA",X"30",X"FA",X"30",X"FA",X"30",X"FA",X"30",X"FA",X"30",X"FA",
		X"30",X"EC",X"2F",X"FA",X"30",X"FA",X"30",X"F9",X"2F",X"FA",X"30",X"FA",X"30",X"FA",X"30",X"FA",
		X"30",X"0A",X"30",X"FA",X"30",X"FA",X"30",X"10",X"09",X"98",X"97",X"10",X"09",X"80",X"A7",X"10",
		X"09",X"28",X"8F",X"13",X"09",X"10",X"8F",X"13",X"08",X"F8",X"AF",X"13",X"08",X"C8",X"9F",X"14",
		X"08",X"50",X"9F",X"11",X"08",X"14",X"AD",X"11",X"08",X"02",X"A7",X"11",X"07",X"F0",X"A3",X"11",
		X"07",X"DE",X"9A",X"11",X"07",X"CC",X"97",X"11",X"07",X"BA",X"90",X"11",X"07",X"78",X"8F",X"11",
		X"07",X"58",X"8F",X"13",X"07",X"40",X"8F",X"10",X"06",X"E0",X"87",X"13",X"06",X"C8",X"87",X"13",
		X"06",X"A0",X"97",X"10",X"06",X"50",X"A7",X"10",X"05",X"60",X"87",X"13",X"05",X"48",X"87",X"13",
		X"05",X"18",X"A7",X"13",X"04",X"B0",X"97",X"14",X"04",X"88",X"9F",X"11",X"04",X"58",X"B3",X"11",
		X"04",X"46",X"AA",X"11",X"04",X"34",X"A7",X"11",X"04",X"22",X"A0",X"11",X"04",X"10",X"97",X"11",
		X"03",X"B8",X"8F",X"13",X"03",X"A0",X"8F",X"13",X"03",X"58",X"9F",X"10",X"02",X"B8",X"8F",X"13",
		X"02",X"A0",X"8F",X"10",X"02",X"88",X"9F",X"13",X"02",X"70",X"9F",X"13",X"01",X"F8",X"97",X"14",
		X"01",X"D0",X"9F",X"11",X"01",X"9C",X"A9",X"11",X"01",X"8A",X"A7",X"11",X"01",X"78",X"9F",X"11",
		X"01",X"66",X"97",X"11",X"01",X"54",X"95",X"11",X"01",X"42",X"8C",X"11",X"00",X"F8",X"AF",X"11",
		X"00",X"E0",X"B7",X"13",X"00",X"B0",X"9F",X"13",X"00",X"48",X"AF",X"FF",X"0D",X"01",X"F0",X"5F",
		X"0D",X"01",X"08",X"67",X"0D",X"00",X"80",X"6F",X"FF",X"0D",X"02",X"30",X"5F",X"0D",X"01",X"80",
		X"5F",X"0D",X"00",X"E8",X"5F",X"0D",X"00",X"18",X"4F",X"FF",X"10",X"09",X"98",X"77",X"13",X"09",
		X"80",X"77",X"10",X"09",X"60",X"7F",X"13",X"09",X"48",X"7F",X"10",X"08",X"E0",X"97",X"10",X"08",
		X"D0",X"7F",X"13",X"08",X"B8",X"7F",X"10",X"08",X"70",X"6F",X"13",X"08",X"58",X"6F",X"13",X"08",
		X"08",X"8F",X"10",X"07",X"E8",X"AF",X"10",X"07",X"C8",X"6F",X"13",X"07",X"B0",X"6F",X"10",X"07",
		X"50",X"97",X"10",X"07",X"40",X"77",X"10",X"07",X"08",X"A7",X"10",X"06",X"E0",X"AF",X"10",X"06",
		X"C8",X"9F",X"10",X"06",X"B0",X"8F",X"10",X"06",X"98",X"87",X"10",X"06",X"78",X"77",X"10",X"06",
		X"48",X"77",X"13",X"06",X"30",X"77",X"10",X"06",X"10",X"67",X"13",X"05",X"F8",X"67",X"13",X"05",
		X"D0",X"B7",X"10",X"05",X"98",X"9F",X"10",X"05",X"88",X"87",X"10",X"05",X"38",X"77",X"13",X"05",
		X"20",X"77",X"10",X"04",X"D8",X"6F",X"13",X"04",X"C0",X"6F",X"10",X"04",X"90",X"77",X"13",X"04",
		X"78",X"77",X"10",X"04",X"38",X"B7",X"10",X"04",X"00",X"77",X"13",X"03",X"E8",X"77",X"10",X"03",
		X"B0",X"97",X"10",X"03",X"90",X"87",X"10",X"03",X"60",X"8F",X"10",X"03",X"30",X"77",X"13",X"03",
		X"18",X"77",X"10",X"02",X"D0",X"7F",X"13",X"02",X"B8",X"7F",X"10",X"02",X"90",X"97",X"10",X"02",
		X"68",X"6F",X"13",X"02",X"50",X"6F",X"10",X"02",X"18",X"8F",X"10",X"01",X"C8",X"77",X"13",X"01",
		X"B0",X"77",X"10",X"01",X"90",X"8F",X"10",X"01",X"58",X"9F",X"10",X"01",X"40",X"6F",X"10",X"01",
		X"10",X"AF",X"10",X"00",X"E0",X"9F",X"10",X"00",X"B8",X"67",X"13",X"00",X"A0",X"67",X"10",X"00",
		X"70",X"87",X"10",X"00",X"48",X"6F",X"13",X"00",X"30",X"6F",X"FF",X"03",X"02",X"00",X"00",X"00",
		X"00",X"00",X"00",X"FD",X"CB",X"24",X"7E",X"28",X"21",X"CD",X"3C",X"31",X"7E",X"FE",X"FF",X"28",
		X"0B",X"CD",X"68",X"31",X"CD",X"8A",X"31",X"FD",X"34",X"6E",X"18",X"ED",X"FD",X"CB",X"24",X"BE",
		X"FD",X"7E",X"28",X"FD",X"77",X"6D",X"FD",X"36",X"6E",X"00",X"CD",X"3C",X"31",X"7E",X"FE",X"FF",
		X"C8",X"CD",X"56",X"31",X"D8",X"CD",X"8A",X"31",X"FD",X"34",X"6E",X"C9",X"FD",X"7E",X"6D",X"E6",
		X"1F",X"87",X"5F",X"16",X"00",X"21",X"F0",X"31",X"19",X"5E",X"23",X"56",X"FD",X"7E",X"6E",X"87",
		X"87",X"6F",X"26",X"00",X"19",X"C9",X"E5",X"23",X"56",X"23",X"5E",X"EB",X"FD",X"56",X"2A",X"FD",
		X"5E",X"2B",X"A7",X"ED",X"52",X"EB",X"E1",X"C9",X"CD",X"56",X"31",X"E5",X"D5",X"FD",X"7E",X"28",
		X"E6",X"0F",X"87",X"5F",X"16",X"00",X"21",X"82",X"1B",X"19",X"5E",X"23",X"56",X"EB",X"56",X"23",
		X"5E",X"EB",X"29",X"29",X"29",X"D1",X"19",X"EB",X"E1",X"C9",X"D5",X"DD",X"21",X"FC",X"63",X"11",
		X"0B",X"00",X"06",X"0C",X"DD",X"CB",X"00",X"7E",X"28",X"06",X"DD",X"19",X"10",X"F6",X"D1",X"C9",
		X"D1",X"7E",X"F6",X"80",X"DD",X"77",X"00",X"E5",X"21",X"00",X"01",X"A7",X"ED",X"52",X"E5",X"2A",
		X"8C",X"63",X"55",X"5C",X"2A",X"A0",X"60",X"A7",X"ED",X"52",X"EB",X"E1",X"7C",X"65",X"FD",X"6E",
		X"2C",X"A7",X"ED",X"52",X"DE",X"00",X"DD",X"77",X"02",X"DD",X"74",X"03",X"DD",X"75",X"04",X"E1",
		X"23",X"23",X"23",X"FD",X"7E",X"2D",X"87",X"87",X"87",X"86",X"DD",X"77",X"05",X"DD",X"36",X"06",
		X"00",X"DD",X"36",X"07",X"00",X"DD",X"36",X"08",X"00",X"3E",X"0C",X"90",X"DD",X"77",X"09",X"C9",
		X"16",X"32",X"86",X"32",X"86",X"32",X"86",X"32",X"86",X"32",X"86",X"32",X"86",X"32",X"37",X"32",
		X"86",X"32",X"44",X"32",X"51",X"32",X"86",X"32",X"86",X"32",X"86",X"32",X"86",X"32",X"86",X"32",
		X"62",X"32",X"86",X"32",X"86",X"32",X"06",X"08",X"A8",X"B7",X"06",X"08",X"28",X"B7",X"06",X"05",
		X"B8",X"A7",X"06",X"05",X"70",X"AF",X"06",X"04",X"6C",X"B7",X"06",X"03",X"20",X"B7",X"06",X"01",
		X"B0",X"B3",X"06",X"00",X"90",X"B7",X"FF",X"06",X"01",X"E0",X"B7",X"06",X"01",X"00",X"B7",X"06",
		X"00",X"20",X"B7",X"FF",X"06",X"01",X"28",X"B7",X"06",X"00",X"C0",X"B7",X"06",X"00",X"70",X"B7",
		X"FF",X"06",X"02",X"08",X"B7",X"06",X"01",X"A0",X"B7",X"06",X"00",X"A8",X"A7",X"06",X"00",X"60",
		X"A7",X"FF",X"06",X"09",X"10",X"8F",X"07",X"07",X"68",X"B7",X"06",X"05",X"B8",X"B7",X"06",X"04",
		X"18",X"9F",X"07",X"03",X"38",X"B7",X"06",X"02",X"70",X"B7",X"06",X"01",X"E8",X"B7",X"06",X"01",
		X"68",X"B7",X"07",X"00",X"F8",X"B7",X"FF",X"DD",X"7E",X"04",X"A7",X"28",X"04",X"DD",X"35",X"04",
		X"C9",X"FD",X"7E",X"0B",X"E6",X"70",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"39",X"33",X"3A",
		X"DC",X"60",X"A7",X"28",X"01",X"23",X"19",X"7E",X"DD",X"77",X"04",X"21",X"49",X"33",X"CB",X"3B",
		X"19",X"DD",X"7E",X"05",X"BE",X"D0",X"CD",X"75",X"07",X"E6",X"01",X"20",X"11",X"CD",X"DF",X"32",
		X"30",X"04",X"CD",X"F1",X"32",X"C9",X"CD",X"EB",X"32",X"D0",X"CD",X"F5",X"32",X"C9",X"CD",X"EB",
		X"32",X"30",X"04",X"CD",X"F5",X"32",X"C9",X"CD",X"DF",X"32",X"D0",X"CD",X"F1",X"32",X"C9",X"FD",
		X"7E",X"14",X"FE",X"11",X"D0",X"FD",X"7E",X"1E",X"FE",X"11",X"C9",X"FD",X"7E",X"32",X"FE",X"11",
		X"C9",X"0E",X"FD",X"18",X"02",X"0E",X"04",X"DD",X"21",X"80",X"64",X"11",X"0A",X"00",X"06",X"08",
		X"DD",X"CB",X"00",X"7E",X"28",X"05",X"DD",X"19",X"10",X"F6",X"C9",X"3E",X"08",X"90",X"CB",X"FF",
		X"CB",X"79",X"28",X"02",X"CB",X"EF",X"DD",X"77",X"00",X"DD",X"71",X"02",X"DD",X"36",X"03",X"00",
		X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"80",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",
		X"DD",X"36",X"08",X"00",X"21",X"F3",X"63",X"34",X"C9",X"40",X"20",X"23",X"19",X"1F",X"17",X"1B",
		X"15",X"17",X"13",X"15",X"12",X"12",X"11",X"10",X"10",X"04",X"05",X"05",X"06",X"06",X"07",X"07",
		X"08",X"3A",X"00",X"60",X"CB",X"77",X"C8",X"21",X"D0",X"64",X"CB",X"7E",X"C0",X"FD",X"7E",X"28",
		X"E6",X"1F",X"C8",X"FE",X"04",X"D0",X"36",X"80",X"E5",X"DD",X"E1",X"DD",X"36",X"02",X"01",X"DD",
		X"36",X"03",X"00",X"DD",X"36",X"04",X"00",X"FD",X"7E",X"2D",X"87",X"87",X"87",X"C6",X"B7",X"DD",
		X"77",X"0B",X"47",X"D6",X"10",X"DD",X"77",X"0A",X"4F",X"FD",X"7E",X"28",X"FE",X"01",X"20",X"05",
		X"DD",X"70",X"05",X"18",X"03",X"DD",X"71",X"05",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",
		X"C9",X"FD",X"7E",X"32",X"E6",X"60",X"FE",X"40",X"C0",X"DD",X"7E",X"06",X"A7",X"28",X"04",X"DD",
		X"35",X"06",X"C9",X"FD",X"7E",X"0B",X"E6",X"70",X"0F",X"0F",X"0F",X"5F",X"16",X"00",X"21",X"39",
		X"33",X"3A",X"DC",X"60",X"A7",X"28",X"01",X"23",X"19",X"7E",X"CB",X"2F",X"CB",X"2F",X"DD",X"77",
		X"06",X"21",X"49",X"33",X"CB",X"3B",X"19",X"DD",X"7E",X"0A",X"BE",X"D0",X"DD",X"21",X"80",X"64",
		X"11",X"0A",X"00",X"06",X"08",X"DD",X"CB",X"00",X"7E",X"28",X"05",X"DD",X"19",X"10",X"F6",X"C9",
		X"3E",X"08",X"90",X"F6",X"88",X"DD",X"77",X"00",X"DD",X"36",X"02",X"04",X"DD",X"36",X"03",X"00",
		X"DD",X"36",X"04",X"00",X"DD",X"36",X"05",X"80",X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",
		X"DD",X"36",X"08",X"00",X"21",X"F8",X"63",X"34",X"3E",X"86",X"32",X"86",X"65",X"C9",X"3A",X"00",
		X"60",X"E6",X"40",X"C8",X"FD",X"7E",X"28",X"FE",X"CC",X"20",X"08",X"FD",X"7E",X"2B",X"FE",X"18",
		X"38",X"10",X"C9",X"E6",X"E0",X"FE",X"C0",X"C0",X"DD",X"7E",X"07",X"A7",X"28",X"04",X"DD",X"35",
		X"07",X"C9",X"FD",X"7E",X"0B",X"E6",X"E0",X"07",X"07",X"07",X"5F",X"16",X"00",X"21",X"9D",X"34",
		X"19",X"7E",X"DD",X"77",X"07",X"21",X"A7",X"34",X"19",X"DD",X"7E",X"08",X"BE",X"D0",X"DD",X"21",
		X"DC",X"64",X"11",X"08",X"00",X"06",X"08",X"DD",X"CB",X"00",X"7E",X"28",X"05",X"DD",X"19",X"10",
		X"F6",X"C9",X"3E",X"08",X"90",X"F6",X"80",X"DD",X"77",X"00",X"DD",X"36",X"02",X"00",X"DD",X"36",
		X"03",X"FF",X"DD",X"36",X"04",X"00",X"CD",X"75",X"07",X"E6",X"0F",X"C6",X"7C",X"DD",X"77",X"05",
		X"DD",X"36",X"06",X"00",X"DD",X"36",X"07",X"00",X"21",X"F6",X"63",X"34",X"C9",X"0D",X"0A",X"09",
		X"09",X"08",X"07",X"07",X"06",X"05",X"05",X"04",X"05",X"05",X"06",X"06",X"07",X"07",X"08",X"08",
		X"08",X"3A",X"00",X"60",X"E6",X"40",X"C8",X"FD",X"7E",X"1E",X"FE",X"49",X"20",X"1E",X"CD",X"24",
		X"35",X"CD",X"33",X"35",X"D0",X"CD",X"75",X"07",X"FD",X"7E",X"20",X"A7",X"20",X"0A",X"FD",X"7E",
		X"21",X"BC",X"30",X"04",X"CB",X"3C",X"BC",X"D8",X"CD",X"61",X"35",X"C9",X"FD",X"7E",X"28",X"FE",
		X"49",X"28",X"0F",X"DD",X"CB",X"00",X"46",X"C8",X"DD",X"CB",X"00",X"86",X"1E",X"15",X"CD",X"0E",
		X"07",X"C9",X"CD",X"24",X"35",X"CD",X"33",X"35",X"D0",X"21",X"C0",X"01",X"FD",X"56",X"2A",X"FD",
		X"5E",X"2B",X"A7",X"ED",X"52",X"EB",X"21",X"00",X"01",X"A7",X"ED",X"52",X"30",X"05",X"CD",X"75",
		X"07",X"18",X"0D",X"7D",X"F5",X"CD",X"75",X"07",X"F1",X"BC",X"38",X"04",X"CB",X"24",X"BC",X"D0",
		X"CD",X"61",X"35",X"C9",X"DD",X"CB",X"00",X"46",X"C0",X"DD",X"CB",X"00",X"C6",X"1E",X"15",X"CD",
		X"FB",X"06",X"C9",X"3A",X"DC",X"60",X"2F",X"E6",X"03",X"28",X"0A",X"DD",X"7E",X"07",X"A7",X"28",
		X"04",X"DD",X"35",X"07",X"C9",X"FD",X"7E",X"0B",X"E6",X"E0",X"07",X"07",X"07",X"5F",X"16",X"00",
		X"21",X"9F",X"34",X"19",X"7E",X"DD",X"77",X"07",X"21",X"A9",X"34",X"19",X"DD",X"7E",X"08",X"BE",
		X"C9",X"DD",X"21",X"DC",X"64",X"11",X"08",X"00",X"06",X"08",X"DD",X"CB",X"00",X"7E",X"28",X"05",
		X"DD",X"19",X"10",X"F6",X"C9",X"DD",X"36",X"02",X"00",X"DD",X"74",X"03",X"DD",X"36",X"04",X"00",
		X"3E",X"08",X"90",X"F6",X"88",X"DD",X"77",X"00",X"DD",X"36",X"05",X"40",X"DD",X"36",X"06",X"00",
		X"DD",X"36",X"07",X"00",X"21",X"F6",X"63",X"34",X"C9",X"45",X"3A",X"54",X"63",X"17",X"D2",X"FE",
		X"35",X"DD",X"CB",X"00",X"6E",X"20",X"23",X"DD",X"CB",X"00",X"EE",X"DD",X"36",X"02",X"00",X"FD",
		X"E5",X"11",X"6F",X"00",X"FD",X"19",X"11",X"08",X"00",X"06",X"18",X"2A",X"A0",X"60",X"FD",X"74",
		X"06",X"FD",X"75",X"07",X"FD",X"19",X"10",X"F6",X"FD",X"E1",X"DD",X"7E",X"02",X"87",X"87",X"87",
		X"5F",X"16",X"00",X"21",X"6F",X"00",X"19",X"EB",X"FD",X"19",X"11",X"18",X"00",X"06",X"03",X"FD",
		X"CB",X"00",X"7E",X"28",X"07",X"D5",X"C5",X"CD",X"1E",X"36",X"C1",X"D1",X"FD",X"19",X"10",X"EF",
		X"DD",X"34",X"02",X"DD",X"7E",X"02",X"FE",X"08",X"D8",X"DD",X"36",X"02",X"00",X"C9",X"11",X"6F",
		X"00",X"FD",X"19",X"11",X"08",X"00",X"06",X"18",X"FD",X"CB",X"00",X"7E",X"28",X"07",X"C5",X"D5",
		X"CD",X"98",X"36",X"D1",X"C1",X"FD",X"19",X"10",X"EF",X"DD",X"36",X"00",X"00",X"C9",X"2A",X"A0",
		X"60",X"FD",X"56",X"06",X"FD",X"5E",X"07",X"FD",X"74",X"06",X"FD",X"75",X"07",X"A7",X"ED",X"52",
		X"EB",X"FD",X"66",X"02",X"FD",X"6E",X"03",X"A7",X"ED",X"52",X"FD",X"74",X"02",X"FD",X"75",X"03",
		X"30",X"04",X"FD",X"35",X"01",X"C9",X"6C",X"FD",X"66",X"01",X"11",X"E0",X"FE",X"19",X"D8",X"FD",
		X"7E",X"00",X"E6",X"07",X"FE",X"01",X"20",X"0F",X"21",X"8A",X"63",X"CB",X"5E",X"20",X"05",X"FD",
		X"35",X"00",X"18",X"03",X"FD",X"34",X"00",X"21",X"FC",X"63",X"11",X"0B",X"00",X"06",X"0C",X"CB",
		X"7E",X"28",X"05",X"19",X"10",X"F9",X"18",X"1B",X"FD",X"7E",X"00",X"77",X"3E",X"0C",X"90",X"EB",
		X"13",X"13",X"FD",X"E5",X"E1",X"23",X"01",X"05",X"00",X"ED",X"B0",X"EB",X"36",X"00",X"23",X"36",
		X"00",X"23",X"77",X"FD",X"36",X"00",X"00",X"C9",X"3A",X"93",X"63",X"67",X"2E",X"00",X"FD",X"56",
		X"06",X"FD",X"5E",X"07",X"A7",X"ED",X"52",X"EB",X"FD",X"66",X"02",X"FD",X"6E",X"03",X"A7",X"ED",
		X"52",X"FD",X"74",X"02",X"FD",X"75",X"03",X"30",X"09",X"CB",X"7A",X"20",X"0C",X"FD",X"35",X"01",
		X"18",X"07",X"CB",X"7A",X"28",X"03",X"FD",X"34",X"01",X"6C",X"FD",X"66",X"01",X"11",X"E0",X"FE",
		X"19",X"D8",X"FD",X"36",X"00",X"00",X"C9",X"3A",X"00",X"60",X"E6",X"40",X"20",X"07",X"3A",X"54",
		X"63",X"17",X"DA",X"37",X"3A",X"CD",X"7B",X"0B",X"30",X"08",X"DD",X"7E",X"02",X"CB",X"7F",X"C2",
		X"37",X"3A",X"DD",X"7E",X"00",X"E6",X"07",X"FE",X"04",X"20",X"34",X"3A",X"8A",X"63",X"E6",X"0C",
		X"20",X"5F",X"DD",X"66",X"02",X"DD",X"6E",X"03",X"11",X"FC",X"FE",X"19",X"38",X"53",X"21",X"8A",
		X"63",X"CB",X"D6",X"21",X"90",X"63",X"36",X"00",X"23",X"DD",X"7E",X"05",X"E6",X"F8",X"0F",X"0F",
		X"0F",X"D6",X"02",X"77",X"23",X"C6",X"02",X"77",X"3E",X"82",X"32",X"86",X"65",X"18",X"32",X"DD",
		X"CB",X"00",X"66",X"C2",X"8C",X"39",X"3A",X"03",X"60",X"DD",X"AE",X"09",X"E6",X"03",X"20",X"48",
		X"DD",X"7E",X"02",X"A7",X"20",X"1B",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"12",X"06",
		X"0F",X"0E",X"0B",X"CD",X"41",X"0A",X"30",X"09",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",X"00",X"E6",
		X"C9",X"DD",X"7E",X"00",X"E6",X"07",X"87",X"5F",X"16",X"00",X"21",X"77",X"37",X"19",X"5E",X"23",
		X"56",X"EB",X"11",X"88",X"37",X"D5",X"E9",X"AD",X"37",X"37",X"3A",X"45",X"38",X"A6",X"38",X"87",
		X"37",X"0F",X"39",X"87",X"37",X"79",X"39",X"C9",X"DD",X"7E",X"02",X"A7",X"C0",X"DD",X"7E",X"00",
		X"E6",X"07",X"87",X"5F",X"16",X"00",X"21",X"C8",X"3A",X"19",X"DD",X"7E",X"07",X"A7",X"28",X"01",
		X"23",X"4E",X"21",X"B8",X"3A",X"19",X"46",X"23",X"56",X"CD",X"02",X"06",X"C9",X"DD",X"7E",X"02",
		X"A7",X"C0",X"DD",X"7E",X"07",X"A7",X"28",X"04",X"DD",X"35",X"07",X"C9",X"FD",X"21",X"54",X"63",
		X"CD",X"15",X"0A",X"C8",X"DD",X"CB",X"00",X"5E",X"20",X"0C",X"DD",X"7E",X"03",X"FE",X"F0",X"D0",
		X"FD",X"BE",X"03",X"D8",X"18",X"32",X"DD",X"7E",X"03",X"FD",X"96",X"03",X"D8",X"C8",X"57",X"ED",
		X"4B",X"E3",X"60",X"CD",X"3C",X"3A",X"7C",X"B5",X"28",X"1E",X"DD",X"7E",X"05",X"FD",X"96",X"05",
		X"D8",X"E5",X"57",X"ED",X"4B",X"7C",X"60",X"CD",X"3C",X"3A",X"EB",X"E1",X"7A",X"B3",X"C8",X"ED",
		X"52",X"38",X"05",X"11",X"F0",X"FF",X"19",X"D8",X"CD",X"CB",X"42",X"C0",X"3E",X"08",X"90",X"F6",
		X"80",X"77",X"E5",X"FD",X"E1",X"FD",X"36",X"02",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"DD",
		X"7E",X"04",X"FD",X"77",X"04",X"DD",X"7E",X"05",X"FD",X"77",X"05",X"FD",X"36",X"06",X"00",X"DD",
		X"7E",X"09",X"FD",X"77",X"07",X"FD",X"36",X"08",X"00",X"3A",X"E1",X"60",X"DD",X"77",X"07",X"1E",
		X"0D",X"CD",X"FB",X"06",X"C9",X"DD",X"7E",X"02",X"A7",X"C0",X"DD",X"7E",X"07",X"A7",X"28",X"04",
		X"DD",X"35",X"07",X"C9",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"C8",X"DD",X"7E",X"03",X"FE",
		X"F0",X"D0",X"FD",X"BE",X"03",X"D8",X"CD",X"CB",X"42",X"C0",X"3E",X"08",X"90",X"F6",X"80",X"77",
		X"E5",X"FD",X"E1",X"FD",X"36",X"02",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"DD",X"7E",X"04",
		X"FD",X"77",X"04",X"DD",X"7E",X"05",X"D6",X"08",X"FD",X"77",X"05",X"FD",X"36",X"06",X"00",X"DD",
		X"7E",X"09",X"F6",X"10",X"FD",X"77",X"07",X"FD",X"36",X"08",X"00",X"FD",X"36",X"09",X"00",X"3A",
		X"E1",X"60",X"DD",X"77",X"07",X"C9",X"3A",X"DC",X"60",X"E6",X"02",X"20",X"05",X"DD",X"CB",X"00",
		X"5E",X"C8",X"DD",X"7E",X"02",X"A7",X"C0",X"DD",X"7E",X"07",X"A7",X"C0",X"FD",X"21",X"54",X"63",
		X"CD",X"15",X"0A",X"C8",X"FD",X"7E",X"03",X"DD",X"96",X"03",X"D8",X"D6",X"10",X"D8",X"CD",X"CB",
		X"42",X"C0",X"3E",X"08",X"90",X"F6",X"80",X"77",X"E5",X"FD",X"E1",X"FD",X"36",X"02",X"00",X"DD",
		X"7E",X"03",X"C6",X"08",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"DD",X"7E",X"05",
		X"D6",X"08",X"FD",X"77",X"05",X"FD",X"36",X"06",X"00",X"DD",X"7E",X"09",X"F6",X"20",X"FD",X"77",
		X"07",X"FD",X"36",X"08",X"00",X"DD",X"36",X"07",X"3C",X"1E",X"0D",X"CD",X"FB",X"06",X"C9",X"DD",
		X"7E",X"02",X"A7",X"C0",X"DD",X"7E",X"07",X"A7",X"28",X"04",X"DD",X"35",X"07",X"C9",X"FD",X"21",
		X"54",X"63",X"CD",X"15",X"0A",X"C8",X"DD",X"7E",X"03",X"FE",X"F0",X"D0",X"FD",X"BE",X"03",X"D8",
		X"CD",X"CB",X"42",X"C0",X"3E",X"08",X"90",X"F6",X"80",X"77",X"E5",X"FD",X"E1",X"FD",X"36",X"02",
		X"00",X"DD",X"7E",X"03",X"D6",X"08",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"DD",
		X"7E",X"05",X"C6",X"08",X"FD",X"77",X"05",X"FD",X"36",X"06",X"00",X"DD",X"7E",X"09",X"F6",X"30",
		X"FD",X"77",X"07",X"FD",X"36",X"08",X"00",X"3A",X"59",X"63",X"FD",X"77",X"09",X"3A",X"E1",X"60",
		X"DD",X"77",X"07",X"1E",X"0D",X"CD",X"FB",X"06",X"C9",X"DD",X"34",X"0A",X"DD",X"CB",X"0A",X"46",
		X"20",X"05",X"DD",X"36",X"07",X"00",X"C9",X"DD",X"36",X"07",X"FF",X"C9",X"DD",X"7E",X"08",X"FE",
		X"0C",X"D2",X"37",X"3A",X"A7",X"20",X"21",X"DD",X"7E",X"00",X"E6",X"07",X"5F",X"87",X"83",X"5F",
		X"16",X"00",X"21",X"DA",X"3A",X"DD",X"7E",X"07",X"A7",X"28",X"03",X"21",X"F2",X"3A",X"19",X"EB",
		X"CD",X"21",X"07",X"1E",X"01",X"CD",X"FB",X"06",X"DD",X"7E",X"08",X"DD",X"34",X"08",X"E6",X"0C",
		X"28",X"06",X"FE",X"04",X"28",X"1B",X"18",X"52",X"01",X"98",X"C0",X"16",X"0D",X"CD",X"02",X"06",
		X"DD",X"7E",X"00",X"E6",X"07",X"FE",X"07",X"C0",X"DD",X"7E",X"08",X"FE",X"02",X"CC",X"56",X"3A",
		X"C9",X"11",X"F8",X"F8",X"CD",X"EF",X"0B",X"01",X"9C",X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",
		X"F8",X"08",X"CD",X"EF",X"0B",X"01",X"A0",X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",X"08",X"F8",
		X"CD",X"EF",X"0B",X"01",X"A4",X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",X"08",X"08",X"CD",X"EF",
		X"0B",X"01",X"EC",X"C0",X"16",X"00",X"CD",X"08",X"06",X"C9",X"11",X"00",X"F8",X"CD",X"EF",X"0B",
		X"01",X"F0",X"C0",X"16",X"02",X"CD",X"08",X"06",X"11",X"00",X"08",X"CD",X"EF",X"0B",X"01",X"F4",
		X"C0",X"16",X"02",X"CD",X"08",X"06",X"C9",X"DD",X"36",X"00",X"00",X"C9",X"3E",X"08",X"1E",X"00",
		X"21",X"00",X"00",X"CB",X"22",X"30",X"04",X"09",X"30",X"01",X"1C",X"3D",X"28",X"05",X"29",X"CB",
		X"13",X"18",X"F0",X"6C",X"63",X"C9",X"11",X"95",X"68",X"21",X"E0",X"D4",X"01",X"40",X"02",X"7E",
		X"12",X"E6",X"08",X"77",X"13",X"23",X"0B",X"78",X"B1",X"20",X"F4",X"1E",X"07",X"CD",X"FB",X"06",
		X"F7",X"CD",X"8B",X"50",X"FD",X"21",X"80",X"64",X"11",X"0A",X"00",X"06",X"08",X"CD",X"15",X"0A",
		X"28",X"0A",X"FD",X"7E",X"02",X"A7",X"20",X"04",X"FD",X"CB",X"00",X"E6",X"FD",X"19",X"10",X"ED",
		X"FD",X"21",X"FC",X"63",X"11",X"0B",X"00",X"06",X"0C",X"CD",X"15",X"0A",X"28",X"0A",X"FD",X"7E",
		X"02",X"A7",X"20",X"04",X"FD",X"CB",X"00",X"E6",X"FD",X"19",X"10",X"ED",X"21",X"95",X"68",X"11",
		X"E0",X"D4",X"01",X"40",X"02",X"ED",X"B0",X"C9",X"C0",X"08",X"80",X"00",X"C0",X"02",X"C0",X"0D",
		X"C0",X"0B",X"F0",X"0D",X"C0",X"00",X"C0",X"00",X"08",X"0C",X"00",X"00",X"30",X"30",X"20",X"24",
		X"48",X"48",X"20",X"24",X"4C",X"4C",X"F8",X"FC",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",
		X"50",X"00",X"00",X"80",X"00",X"00",X"00",X"00",X"00",X"80",X"00",X"01",X"00",X"00",X"03",X"00",
		X"00",X"00",X"50",X"00",X"00",X"00",X"00",X"00",X"50",X"00",X"00",X"50",X"00",X"00",X"00",X"00",
		X"00",X"50",X"00",X"01",X"00",X"00",X"03",X"00",X"DD",X"CB",X"00",X"5E",X"C2",X"BA",X"3E",X"DD",
		X"7E",X"02",X"A7",X"28",X"07",X"3A",X"54",X"63",X"17",X"D2",X"52",X"3E",X"DD",X"CB",X"00",X"66",
		X"C2",X"A6",X"3D",X"06",X"05",X"CD",X"7A",X"06",X"DD",X"7E",X"02",X"A7",X"28",X"62",X"FA",X"19",
		X"3D",X"DD",X"CB",X"00",X"6E",X"20",X"1F",X"CD",X"7B",X"0B",X"FD",X"7E",X"28",X"FE",X"11",X"DC",
		X"85",X"0B",X"FD",X"7E",X"28",X"FD",X"46",X"2D",X"CD",X"5B",X"3E",X"DD",X"7E",X"02",X"A7",X"C0",
		X"1E",X"10",X"CD",X"FB",X"06",X"C9",X"FD",X"7E",X"32",X"FE",X"11",X"30",X"29",X"21",X"00",X"08",
		X"ED",X"5B",X"7C",X"60",X"A7",X"ED",X"52",X"DD",X"56",X"03",X"DD",X"5E",X"04",X"19",X"DD",X"74",
		X"03",X"DD",X"75",X"04",X"30",X"0A",X"DD",X"34",X"02",X"DD",X"7E",X"02",X"FE",X"02",X"30",X"06",
		X"06",X"80",X"CD",X"6A",X"3E",X"C9",X"DD",X"CB",X"00",X"AE",X"3E",X"80",X"32",X"86",X"65",X"C9",
		X"DD",X"CB",X"00",X"6E",X"28",X"31",X"FD",X"7E",X"28",X"FE",X"11",X"30",X"26",X"ED",X"5B",X"7C",
		X"60",X"CB",X"3A",X"CB",X"1B",X"21",X"00",X"04",X"A7",X"ED",X"52",X"DD",X"56",X"03",X"DD",X"5E",
		X"04",X"19",X"DD",X"74",X"03",X"DD",X"75",X"04",X"30",X"36",X"DD",X"34",X"02",X"1E",X"10",X"CD",
		X"0E",X"07",X"C9",X"DD",X"CB",X"00",X"AE",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"ED",X"5B",X"7C",
		X"60",X"7A",X"B3",X"20",X"05",X"11",X"00",X"04",X"18",X"0B",X"FD",X"7E",X"1E",X"FE",X"11",X"38",
		X"04",X"CB",X"3A",X"CB",X"1B",X"CD",X"85",X"0B",X"30",X"06",X"1E",X"10",X"CD",X"0E",X"07",X"C9",
		X"FD",X"7E",X"20",X"A7",X"20",X"08",X"FD",X"7E",X"21",X"DD",X"BE",X"03",X"38",X"0B",X"FD",X"7E",
		X"1E",X"FD",X"46",X"23",X"CD",X"5B",X"3E",X"18",X"09",X"FD",X"7E",X"28",X"FD",X"46",X"2D",X"CD",
		X"5B",X"3E",X"06",X"C0",X"0E",X"04",X"16",X"01",X"CD",X"02",X"06",X"3A",X"03",X"60",X"DD",X"AE",
		X"00",X"E6",X"03",X"C0",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",X"0A",X"06",X"0F",X"0E",
		X"07",X"CD",X"41",X"0A",X"DA",X"BA",X"3C",X"FD",X"21",X"60",X"63",X"CD",X"15",X"0A",X"28",X"09",
		X"06",X"18",X"0E",X"05",X"CD",X"41",X"0A",X"38",X"71",X"FD",X"21",X"68",X"63",X"CD",X"15",X"0A",
		X"28",X"0F",X"FD",X"CB",X"00",X"46",X"20",X"09",X"06",X"0B",X"0E",X"05",X"CD",X"41",X"0A",X"38",
		X"59",X"FD",X"21",X"79",X"63",X"CD",X"15",X"0A",X"28",X"0F",X"FD",X"CB",X"00",X"46",X"20",X"09",
		X"06",X"0B",X"0E",X"05",X"CD",X"41",X"0A",X"38",X"41",X"FD",X"21",X"D0",X"64",X"CD",X"15",X"0A",
		X"28",X"09",X"06",X"0F",X"0E",X"0A",X"CD",X"41",X"0A",X"38",X"2F",X"DD",X"7E",X"00",X"E6",X"07",
		X"28",X"31",X"FD",X"21",X"BC",X"64",X"11",X"F6",X"FF",X"67",X"D6",X"07",X"28",X"07",X"ED",X"44",
		X"FD",X"19",X"3D",X"20",X"FB",X"06",X"10",X"0E",X"08",X"CD",X"15",X"0A",X"28",X"05",X"CD",X"41",
		X"0A",X"38",X"07",X"FD",X"19",X"25",X"20",X"F1",X"18",X"09",X"FD",X"CB",X"00",X"E6",X"DD",X"CB",
		X"00",X"E6",X"C9",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"C8",X"DD",X"7E",X"08",X"A7",X"28",
		X"04",X"DD",X"35",X"08",X"C9",X"CD",X"CB",X"42",X"C0",X"3E",X"08",X"90",X"F6",X"80",X"77",X"E5",
		X"FD",X"E1",X"FD",X"36",X"02",X"00",X"DD",X"7E",X"03",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",
		X"77",X"04",X"DD",X"7E",X"05",X"FD",X"77",X"05",X"DD",X"7E",X"06",X"FD",X"77",X"06",X"DD",X"7E",
		X"00",X"E6",X"07",X"F6",X"40",X"FD",X"77",X"07",X"FD",X"36",X"08",X"00",X"CD",X"DA",X"42",X"DD",
		X"36",X"08",X"08",X"1E",X"0F",X"CD",X"FB",X"06",X"C9",X"DD",X"CB",X"00",X"6E",X"20",X"30",X"CD",
		X"7B",X"0B",X"FD",X"7E",X"14",X"FE",X"11",X"DC",X"85",X"0B",X"06",X"80",X"CD",X"6A",X"3E",X"DD",
		X"7E",X"02",X"FE",X"FF",X"D0",X"FE",X"FD",X"DA",X"52",X"3E",X"FD",X"7E",X"1E",X"FE",X"11",X"D0",
		X"DD",X"CB",X"00",X"EE",X"1E",X"0C",X"CD",X"FB",X"06",X"3E",X"80",X"32",X"86",X"65",X"C9",X"FD",
		X"7E",X"1E",X"FE",X"11",X"30",X"46",X"21",X"00",X"08",X"ED",X"5B",X"7C",X"60",X"A7",X"ED",X"52",
		X"DD",X"56",X"03",X"DD",X"5E",X"04",X"19",X"DD",X"74",X"03",X"DD",X"75",X"04",X"30",X"23",X"DD",
		X"34",X"02",X"DD",X"7E",X"02",X"A7",X"28",X"10",X"FE",X"FE",X"20",X"16",X"1E",X"0C",X"CD",X"FB",
		X"06",X"3E",X"80",X"32",X"86",X"65",X"18",X"0A",X"1E",X"10",X"CD",X"FB",X"06",X"1E",X"0C",X"CD",
		X"0E",X"07",X"FD",X"7E",X"1E",X"FD",X"46",X"23",X"CD",X"5B",X"3E",X"C9",X"DD",X"CB",X"00",X"AE",
		X"1E",X"0C",X"CD",X"0E",X"07",X"C9",X"DD",X"7E",X"07",X"FE",X"0C",X"D2",X"52",X"3E",X"A7",X"20",
		X"10",X"11",X"92",X"40",X"CD",X"21",X"07",X"1E",X"10",X"CD",X"0E",X"07",X"1E",X"0A",X"CD",X"FB",
		X"06",X"CD",X"7B",X"0B",X"DA",X"52",X"3E",X"DD",X"7E",X"07",X"DD",X"34",X"07",X"E6",X"0C",X"28",
		X"06",X"FE",X"04",X"28",X"0B",X"18",X"42",X"01",X"A8",X"C0",X"16",X"0F",X"CD",X"02",X"06",X"C9",
		X"11",X"F8",X"F8",X"CD",X"EF",X"0B",X"01",X"AC",X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",X"F8",
		X"08",X"CD",X"EF",X"0B",X"01",X"B0",X"C0",X"16",X"00",X"CD",X"08",X"06",X"11",X"08",X"F8",X"CD",
		X"EF",X"0B",X"01",X"B0",X"F0",X"16",X"00",X"CD",X"08",X"06",X"11",X"08",X"08",X"CD",X"EF",X"0B",
		X"01",X"AC",X"F0",X"16",X"00",X"CD",X"08",X"06",X"C9",X"11",X"F8",X"F8",X"CD",X"EF",X"0B",X"01",
		X"B4",X"C0",X"16",X"0C",X"CD",X"08",X"06",X"11",X"F8",X"08",X"CD",X"EF",X"0B",X"01",X"B8",X"C0",
		X"16",X"0C",X"CD",X"08",X"06",X"11",X"08",X"F8",X"CD",X"EF",X"0B",X"01",X"B8",X"F0",X"16",X"0C",
		X"CD",X"08",X"06",X"11",X"08",X"08",X"CD",X"EF",X"0B",X"01",X"B4",X"F0",X"16",X"0C",X"CD",X"08",
		X"06",X"C9",X"DD",X"36",X"00",X"00",X"21",X"F3",X"63",X"35",X"C9",X"E6",X"1F",X"5F",X"16",X"00",
		X"21",X"A7",X"3E",X"19",X"78",X"87",X"87",X"87",X"86",X"47",X"DD",X"34",X"09",X"DD",X"7E",X"05",
		X"FE",X"40",X"38",X"09",X"B8",X"30",X"1B",X"DD",X"CB",X"09",X"7E",X"20",X"15",X"DD",X"66",X"05",
		X"DD",X"6E",X"06",X"11",X"00",X"01",X"19",X"DD",X"74",X"05",X"DD",X"75",X"06",X"DD",X"CB",X"09",
		X"BE",X"C9",X"DD",X"66",X"05",X"DD",X"6E",X"06",X"11",X"00",X"FF",X"19",X"DD",X"74",X"05",X"DD",
		X"75",X"06",X"DD",X"CB",X"09",X"FE",X"C9",X"70",X"B0",X"A8",X"A8",X"A8",X"70",X"38",X"88",X"38",
		X"88",X"88",X"38",X"78",X"38",X"70",X"38",X"58",X"88",X"38",X"DD",X"7E",X"02",X"A7",X"28",X"07",
		X"3A",X"54",X"63",X"17",X"D2",X"49",X"40",X"DD",X"CB",X"00",X"66",X"C2",X"27",X"40",X"06",X"05",
		X"CD",X"7A",X"06",X"DD",X"7E",X"02",X"A7",X"FA",X"12",X"40",X"28",X"1B",X"CD",X"7B",X"0B",X"FD",
		X"7E",X"28",X"E6",X"60",X"FE",X"40",X"CC",X"85",X"0B",X"CD",X"52",X"40",X"DD",X"7E",X"02",X"A7",
		X"C0",X"1E",X"14",X"CD",X"FB",X"06",X"C9",X"ED",X"5B",X"7C",X"60",X"7A",X"B3",X"20",X"03",X"11",
		X"00",X"04",X"DD",X"66",X"03",X"DD",X"6E",X"04",X"CD",X"85",X"0B",X"30",X"06",X"1E",X"14",X"CD",
		X"0E",X"07",X"C9",X"CD",X"52",X"40",X"06",X"C0",X"0E",X"68",X"16",X"0B",X"CD",X"02",X"06",X"3A",
		X"03",X"60",X"DD",X"AE",X"00",X"E6",X"03",X"C0",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"28",
		X"09",X"06",X"0F",X"0E",X"07",X"CD",X"41",X"0A",X"38",X"71",X"FD",X"21",X"60",X"63",X"CD",X"15",
		X"0A",X"28",X"09",X"06",X"18",X"0E",X"05",X"CD",X"41",X"0A",X"38",X"5F",X"FD",X"21",X"68",X"63",
		X"CD",X"15",X"0A",X"28",X"0F",X"FD",X"CB",X"00",X"46",X"20",X"09",X"06",X"0B",X"0E",X"05",X"CD",
		X"41",X"0A",X"38",X"47",X"FD",X"21",X"79",X"63",X"CD",X"15",X"0A",X"28",X"0F",X"FD",X"CB",X"00",
		X"46",X"20",X"09",X"06",X"0B",X"0E",X"05",X"CD",X"41",X"0A",X"38",X"2F",X"DD",X"7E",X"00",X"E6",
		X"07",X"28",X"31",X"FD",X"21",X"BC",X"64",X"11",X"F6",X"FF",X"67",X"D6",X"07",X"28",X"07",X"ED",
		X"44",X"FD",X"19",X"3D",X"20",X"FB",X"06",X"10",X"0E",X"08",X"CD",X"15",X"0A",X"28",X"05",X"CD",
		X"41",X"0A",X"38",X"07",X"FD",X"19",X"25",X"20",X"F1",X"18",X"09",X"DD",X"CB",X"00",X"E6",X"FD",
		X"CB",X"00",X"E6",X"C9",X"FD",X"21",X"54",X"63",X"CD",X"15",X"0A",X"C8",X"DD",X"7E",X"08",X"A7",
		X"28",X"04",X"DD",X"35",X"08",X"C9",X"3A",X"57",X"63",X"DD",X"BE",X"03",X"D0",X"CD",X"CB",X"42",
		X"C0",X"3E",X"08",X"90",X"F6",X"80",X"77",X"E5",X"FD",X"E1",X"FD",X"36",X"02",X"00",X"DD",X"7E",
		X"03",X"D6",X"08",X"FD",X"77",X"03",X"DD",X"7E",X"04",X"FD",X"77",X"04",X"DD",X"7E",X"05",X"C6",
		X"02",X"FD",X"77",X"05",X"DD",X"7E",X"06",X"FD",X"77",X"06",X"DD",X"7E",X"00",X"E6",X"07",X"F6");
begin
process(clk)
begin
	if rising_edge(clk) then
		data <= rom_data(to_integer(unsigned(addr)));
	end if;
end process;
end architecture;
